module Data_Mem (
MemRead_i, 
MemWrite_i, 
\addr_i[0], 
\addr_i[10], 
\addr_i[11], 
\addr_i[12], 
\addr_i[13], 
\addr_i[14], 
\addr_i[15], 
\addr_i[16], 
\addr_i[17], 
\addr_i[18], 
\addr_i[19], 
\addr_i[1], 
\addr_i[20], 
\addr_i[21], 
\addr_i[22], 
\addr_i[23], 
\addr_i[24], 
\addr_i[25], 
\addr_i[26], 
\addr_i[27], 
\addr_i[28], 
\addr_i[29], 
\addr_i[2], 
\addr_i[30], 
\addr_i[31], 
\addr_i[3], 
\addr_i[4], 
\addr_i[5], 
\addr_i[6], 
\addr_i[7], 
\addr_i[8], 
\addr_i[9], 
\data_i[0], 
\data_i[10], 
\data_i[11], 
\data_i[12], 
\data_i[13], 
\data_i[14], 
\data_i[15], 
\data_i[16], 
\data_i[17], 
\data_i[18], 
\data_i[19], 
\data_i[1], 
\data_i[20], 
\data_i[21], 
\data_i[22], 
\data_i[23], 
\data_i[24], 
\data_i[25], 
\data_i[26], 
\data_i[27], 
\data_i[28], 
\data_i[29], 
\data_i[2], 
\data_i[30], 
\data_i[31], 
\data_i[3], 
\data_i[4], 
\data_i[5], 
\data_i[6], 
\data_i[7], 
\data_i[8], 
\data_i[9], 
\memory[0][0], 
\memory[0][1], 
\memory[0][2], 
\memory[0][3], 
\memory[0][4], 
\memory[0][5], 
\memory[0][6], 
\memory[0][7], 
\memory[10][0], 
\memory[10][1], 
\memory[10][2], 
\memory[10][3], 
\memory[10][4], 
\memory[10][5], 
\memory[10][6], 
\memory[10][7], 
\memory[11][0], 
\memory[11][1], 
\memory[11][2], 
\memory[11][3], 
\memory[11][4], 
\memory[11][5], 
\memory[11][6], 
\memory[11][7], 
\memory[12][0], 
\memory[12][1], 
\memory[12][2], 
\memory[12][3], 
\memory[12][4], 
\memory[12][5], 
\memory[12][6], 
\memory[12][7], 
\memory[13][0], 
\memory[13][1], 
\memory[13][2], 
\memory[13][3], 
\memory[13][4], 
\memory[13][5], 
\memory[13][6], 
\memory[13][7], 
\memory[14][0], 
\memory[14][1], 
\memory[14][2], 
\memory[14][3], 
\memory[14][4], 
\memory[14][5], 
\memory[14][6], 
\memory[14][7], 
\memory[15][0], 
\memory[15][1], 
\memory[15][2], 
\memory[15][3], 
\memory[15][4], 
\memory[15][5], 
\memory[15][6], 
\memory[15][7], 
\memory[16][0], 
\memory[16][1], 
\memory[16][2], 
\memory[16][3], 
\memory[16][4], 
\memory[16][5], 
\memory[16][6], 
\memory[16][7], 
\memory[17][0], 
\memory[17][1], 
\memory[17][2], 
\memory[17][3], 
\memory[17][4], 
\memory[17][5], 
\memory[17][6], 
\memory[17][7], 
\memory[18][0], 
\memory[18][1], 
\memory[18][2], 
\memory[18][3], 
\memory[18][4], 
\memory[18][5], 
\memory[18][6], 
\memory[18][7], 
\memory[19][0], 
\memory[19][1], 
\memory[19][2], 
\memory[19][3], 
\memory[19][4], 
\memory[19][5], 
\memory[19][6], 
\memory[19][7], 
\memory[1][0], 
\memory[1][1], 
\memory[1][2], 
\memory[1][3], 
\memory[1][4], 
\memory[1][5], 
\memory[1][6], 
\memory[1][7], 
\memory[20][0], 
\memory[20][1], 
\memory[20][2], 
\memory[20][3], 
\memory[20][4], 
\memory[20][5], 
\memory[20][6], 
\memory[20][7], 
\memory[21][0], 
\memory[21][1], 
\memory[21][2], 
\memory[21][3], 
\memory[21][4], 
\memory[21][5], 
\memory[21][6], 
\memory[21][7], 
\memory[22][0], 
\memory[22][1], 
\memory[22][2], 
\memory[22][3], 
\memory[22][4], 
\memory[22][5], 
\memory[22][6], 
\memory[22][7], 
\memory[23][0], 
\memory[23][1], 
\memory[23][2], 
\memory[23][3], 
\memory[23][4], 
\memory[23][5], 
\memory[23][6], 
\memory[23][7], 
\memory[24][0], 
\memory[24][1], 
\memory[24][2], 
\memory[24][3], 
\memory[24][4], 
\memory[24][5], 
\memory[24][6], 
\memory[24][7], 
\memory[25][0], 
\memory[25][1], 
\memory[25][2], 
\memory[25][3], 
\memory[25][4], 
\memory[25][5], 
\memory[25][6], 
\memory[25][7], 
\memory[26][0], 
\memory[26][1], 
\memory[26][2], 
\memory[26][3], 
\memory[26][4], 
\memory[26][5], 
\memory[26][6], 
\memory[26][7], 
\memory[27][0], 
\memory[27][1], 
\memory[27][2], 
\memory[27][3], 
\memory[27][4], 
\memory[27][5], 
\memory[27][6], 
\memory[27][7], 
\memory[28][0], 
\memory[28][1], 
\memory[28][2], 
\memory[28][3], 
\memory[28][4], 
\memory[28][5], 
\memory[28][6], 
\memory[28][7], 
\memory[29][0], 
\memory[29][1], 
\memory[29][2], 
\memory[29][3], 
\memory[29][4], 
\memory[29][5], 
\memory[29][6], 
\memory[29][7], 
\memory[2][0], 
\memory[2][1], 
\memory[2][2], 
\memory[2][3], 
\memory[2][4], 
\memory[2][5], 
\memory[2][6], 
\memory[2][7], 
\memory[30][0], 
\memory[30][1], 
\memory[30][2], 
\memory[30][3], 
\memory[30][4], 
\memory[30][5], 
\memory[30][6], 
\memory[30][7], 
\memory[31][0], 
\memory[31][1], 
\memory[31][2], 
\memory[31][3], 
\memory[31][4], 
\memory[31][5], 
\memory[31][6], 
\memory[31][7], 
\memory[3][0], 
\memory[3][1], 
\memory[3][2], 
\memory[3][3], 
\memory[3][4], 
\memory[3][5], 
\memory[3][6], 
\memory[3][7], 
\memory[4][0], 
\memory[4][1], 
\memory[4][2], 
\memory[4][3], 
\memory[4][4], 
\memory[4][5], 
\memory[4][6], 
\memory[4][7], 
\memory[5][0], 
\memory[5][1], 
\memory[5][2], 
\memory[5][3], 
\memory[5][4], 
\memory[5][5], 
\memory[5][6], 
\memory[5][7], 
\memory[6][0], 
\memory[6][1], 
\memory[6][2], 
\memory[6][3], 
\memory[6][4], 
\memory[6][5], 
\memory[6][6], 
\memory[6][7], 
\memory[7][0], 
\memory[7][1], 
\memory[7][2], 
\memory[7][3], 
\memory[7][4], 
\memory[7][5], 
\memory[7][6], 
\memory[7][7], 
\memory[8][0], 
\memory[8][1], 
\memory[8][2], 
\memory[8][3], 
\memory[8][4], 
\memory[8][5], 
\memory[8][6], 
\memory[8][7], 
\memory[9][0], 
\memory[9][1], 
\memory[9][2], 
\memory[9][3], 
\memory[9][4], 
\memory[9][5], 
\memory[9][6], 
\memory[9][7], 
\op_addr[0], 
\op_addr[1], 
\op_addr[2], 
\op_addr[3], 
\op_addr[4], 
clk_i, 
reset,
\data_mem_o[0], 
\data_mem_o[10], 
\data_mem_o[11], 
\data_mem_o[12], 
\data_mem_o[13], 
\data_mem_o[14], 
\data_mem_o[15], 
\data_mem_o[16], 
\data_mem_o[17], 
\data_mem_o[18], 
\data_mem_o[19], 
\data_mem_o[1], 
\data_mem_o[20], 
\data_mem_o[21], 
\data_mem_o[22], 
\data_mem_o[23], 
\data_mem_o[24], 
\data_mem_o[25], 
\data_mem_o[26], 
\data_mem_o[27], 
\data_mem_o[28], 
\data_mem_o[29], 
\data_mem_o[2], 
\data_mem_o[30], 
\data_mem_o[31], 
\data_mem_o[3], 
\data_mem_o[4], 
\data_mem_o[5], 
\data_mem_o[6], 
\data_mem_o[7], 
\data_mem_o[8], 
\data_mem_o[9], 
\data_o[0], 
\data_o[10], 
\data_o[11], 
\data_o[12], 
\data_o[13], 
\data_o[14], 
\data_o[15], 
\data_o[16], 
\data_o[17], 
\data_o[18], 
\data_o[19], 
\data_o[1], 
\data_o[20], 
\data_o[21], 
\data_o[22], 
\data_o[23], 
\data_o[24], 
\data_o[25], 
\data_o[26], 
\data_o[27], 
\data_o[28], 
\data_o[29], 
\data_o[2], 
\data_o[30], 
\data_o[31], 
\data_o[3], 
\data_o[4], 
\data_o[5], 
\data_o[6], 
\data_o[7], 
\data_o[8], 
\data_o[9], 
_00000_, 
_00001_, 
_00002_, 
_00003_, 
_00004_, 
_00005_, 
_00006_, 
_00007_, 
_00008_, 
_00009_, 
_00010_, 
_00011_, 
_00012_, 
_00013_, 
_00014_, 
_00015_, 
_00016_, 
_00017_, 
_00018_, 
_00019_, 
_00020_, 
_00021_, 
_00022_, 
_00023_, 
_00024_, 
_00025_, 
_00026_, 
_00027_, 
_00028_, 
_00029_, 
_00030_, 
_00031_, 
_00032_, 
_00033_, 
_00034_, 
_00035_, 
_00036_, 
_00037_, 
_00038_, 
_00039_, 
_00040_, 
_00041_, 
_00042_, 
_00043_, 
_00044_, 
_00045_, 
_00046_, 
_00047_, 
_00048_, 
_00049_, 
_00050_, 
_00051_, 
_00052_, 
_00053_, 
_00054_, 
_00055_, 
_00056_, 
_00057_, 
_00058_, 
_00059_, 
_00060_, 
_00061_, 
_00062_, 
_00063_, 
_00064_, 
_00065_, 
_00066_, 
_00067_, 
_00068_, 
_00069_, 
_00070_, 
_00071_, 
_00072_, 
_00073_, 
_00074_, 
_00075_, 
_00076_, 
_00077_, 
_00078_, 
_00079_, 
_00080_, 
_00081_, 
_00082_, 
_00083_, 
_00084_, 
_00085_, 
_00086_, 
_00087_, 
_00088_, 
_00089_, 
_00090_, 
_00091_, 
_00092_, 
_00093_, 
_00094_, 
_00095_, 
_00096_, 
_00097_, 
_00098_, 
_00099_, 
_00100_, 
_00101_, 
_00102_, 
_00103_, 
_00104_, 
_00105_, 
_00106_, 
_00107_, 
_00108_, 
_00109_, 
_00110_, 
_00111_, 
_00112_, 
_00113_, 
_00114_, 
_00115_, 
_00116_, 
_00117_, 
_00118_, 
_00119_, 
_00120_, 
_00121_, 
_00122_, 
_00123_, 
_00124_, 
_00125_, 
_00126_, 
_00127_, 
_00128_, 
_00129_, 
_00130_, 
_00131_, 
_00132_, 
_00133_, 
_00134_, 
_00135_, 
_00136_, 
_00137_, 
_00138_, 
_00139_, 
_00140_, 
_00141_, 
_00142_, 
_00143_, 
_00144_, 
_00145_, 
_00146_, 
_00147_, 
_00148_, 
_00149_, 
_00150_, 
_00151_, 
_00152_, 
_00153_, 
_00154_, 
_00155_, 
_00156_, 
_00157_, 
_00158_, 
_00159_, 
_00160_, 
_00161_, 
_00162_, 
_00163_, 
_00164_, 
_00165_, 
_00166_, 
_00167_, 
_00168_, 
_00169_, 
_00170_, 
_00171_, 
_00172_, 
_00173_, 
_00174_, 
_00175_, 
_00176_, 
_00177_, 
_00178_, 
_00179_, 
_00180_, 
_00181_, 
_00182_, 
_00183_, 
_00184_, 
_00185_, 
_00186_, 
_00187_, 
_00188_, 
_00189_, 
_00190_, 
_00191_, 
_00192_, 
_00193_, 
_00194_, 
_00195_, 
_00196_, 
_00197_, 
_00198_, 
_00199_, 
_00200_, 
_00201_, 
_00202_, 
_00203_, 
_00204_, 
_00205_, 
_00206_, 
_00207_, 
_00208_, 
_00209_, 
_00210_, 
_00211_, 
_00212_, 
_00213_, 
_00214_, 
_00215_, 
_00216_, 
_00217_, 
_00218_, 
_00219_, 
_00220_, 
_00221_, 
_00222_, 
_00223_, 
_00224_, 
_00225_, 
_00226_, 
_00227_, 
_00228_, 
_00229_, 
_00230_, 
_00231_, 
_00232_, 
_00233_, 
_00234_, 
_00235_, 
_00236_, 
_00237_, 
_00238_, 
_00239_, 
_00240_, 
_00241_, 
_00242_, 
_00243_, 
_00244_, 
_00245_, 
_00246_, 
_00247_, 
_00248_, 
_00249_, 
_00250_, 
_00251_, 
_00252_, 
_00253_, 
_00254_, 
_00255_
);
  wire _00256_;
  wire _00257_;
  wire _00258_;
  wire _00259_;
  wire _00260_;
  wire _00261_;
  wire _00262_;
  wire _00263_;
  wire _00264_;
  wire _00265_;
  wire _00266_;
  wire _00267_;
  wire _00268_;
  wire _00269_;
  wire _00270_;
  wire _00271_;
  wire _00272_;
  wire _00273_;
  wire _00274_;
  wire _00275_;
  wire _00276_;
  wire _00277_;
  wire _00278_;
  wire _00279_;
  wire _00280_;
  wire _00281_;
  wire _00282_;
  wire _00283_;
  wire _00284_;
  wire _00285_;
  wire _00286_;
  wire _00287_;
  wire _00288_;
  wire _00289_;
  wire _00290_;
  wire _00291_;
  wire _00292_;
  wire _00293_;
  wire _00294_;
  wire _00295_;
  wire _00296_;
  wire _00297_;
  wire _00298_;
  wire _00299_;
  wire _00300_;
  wire _00301_;
  wire _00302_;
  wire _00303_;
  wire _00304_;
  wire _00305_;
  wire _00306_;
  wire _00307_;
  wire _00308_;
  wire _00309_;
  wire _00310_;
  wire _00311_;
  wire _00312_;
  wire _00313_;
  wire _00314_;
  wire _00315_;
  wire _00316_;
  wire _00317_;
  wire _00318_;
  wire _00319_;
  wire _00320_;
  wire _00321_;
  wire _00322_;
  wire _00323_;
  wire _00324_;
  wire _00325_;
  wire _00326_;
  wire _00327_;
  wire _00328_;
  wire _00329_;
  wire _00330_;
  wire _00331_;
  wire _00332_;
  wire _00333_;
  wire _00334_;
  wire _00335_;
  wire _00336_;
  wire _00337_;
  wire _00338_;
  wire _00339_;
  wire _00340_;
  wire _00341_;
  wire _00342_;
  wire _00343_;
  wire _00344_;
  wire _00345_;
  wire _00346_;
  wire _00347_;
  wire _00348_;
  wire _00349_;
  wire _00350_;
  wire _00351_;
  wire _00352_;
  wire _00353_;
  wire _00354_;
  wire _00355_;
  wire _00356_;
  wire _00357_;
  wire _00358_;
  wire _00359_;
  wire _00360_;
  wire _00361_;
  wire _00362_;
  wire _00363_;
  wire _00364_;
  wire _00365_;
  wire _00366_;
  wire _00367_;
  wire _00368_;
  wire _00369_;
  wire _00370_;
  wire _00371_;
  wire _00372_;
  wire _00373_;
  wire _00374_;
  wire _00375_;
  wire _00376_;
  wire _00377_;
  wire _00378_;
  wire _00379_;
  wire _00380_;
  wire _00381_;
  wire _00382_;
  wire _00383_;
  wire _00384_;
  wire _00385_;
  wire _00386_;
  wire _00387_;
  wire _00388_;
  wire _00389_;
  wire _00390_;
  wire _00391_;
  wire _00392_;
  wire _00393_;
  wire _00394_;
  wire _00395_;
  wire _00396_;
  wire _00397_;
  wire _00398_;
  wire _00399_;
  wire _00400_;
  wire _00401_;
  wire _00402_;
  wire _00403_;
  wire _00404_;
  wire _00405_;
  wire _00406_;
  wire _00407_;
  wire _00408_;
  wire _00409_;
  wire _00410_;
  wire _00411_;
  wire _00412_;
  wire _00413_;
  wire _00414_;
  wire _00415_;
  wire _00416_;
  wire _00417_;
  wire _00418_;
  wire _00419_;
  wire _00420_;
  wire _00421_;
  wire _00422_;
  wire _00423_;
  wire _00424_;
  wire _00425_;
  wire _00426_;
  wire _00427_;
  wire _00428_;
  wire _00429_;
  wire _00430_;
  wire _00431_;
  wire _00432_;
  wire _00433_;
  wire _00434_;
  wire _00435_;
  wire _00436_;
  wire _00437_;
  wire _00438_;
  wire _00439_;
  wire _00440_;
  wire _00441_;
  wire _00442_;
  wire _00443_;
  wire _00444_;
  wire _00445_;
  wire _00446_;
  wire _00447_;
  wire _00448_;
  wire _00449_;
  wire _00450_;
  wire _00451_;
  wire _00452_;
  wire _00453_;
  wire _00454_;
  wire _00455_;
  wire _00456_;
  wire _00457_;
  wire _00458_;
  wire _00459_;
  wire _00460_;
  wire _00461_;
  wire _00462_;
  wire _00463_;
  wire _00464_;
  wire _00465_;
  wire _00466_;
  wire _00467_;
  wire _00468_;
  wire _00469_;
  wire _00470_;
  wire _00471_;
  wire _00472_;
  wire _00473_;
  wire _00474_;
  wire _00475_;
  wire _00476_;
  wire _00477_;
  wire _00478_;
  wire _00479_;
  wire _00480_;
  wire _00481_;
  wire _00482_;
  wire _00483_;
  wire _00484_;
  wire _00485_;
  wire _00486_;
  wire _00487_;
  wire _00488_;
  wire _00489_;
  wire _00490_;
  wire _00491_;
  wire _00492_;
  wire _00493_;
  wire _00494_;
  wire _00495_;
  wire _00496_;
  wire _00497_;
  wire _00498_;
  wire _00499_;
  wire _00500_;
  wire _00501_;
  wire _00502_;
  wire _00503_;
  wire _00504_;
  wire _00505_;
  wire _00506_;
  wire _00507_;
  wire _00508_;
  wire _00509_;
  wire _00510_;
  wire _00511_;
  wire _00512_;
  wire _00513_;
  wire _00514_;
  wire _00515_;
  wire _00516_;
  wire _00517_;
  wire _00518_;
  wire _00519_;
  wire _00520_;
  wire _00521_;
  wire _00522_;
  wire _00523_;
  wire _00524_;
  wire _00525_;
  wire _00526_;
  wire _00527_;
  wire _00528_;
  wire _00529_;
  wire _00530_;
  wire _00531_;
  wire _00532_;
  wire _00533_;
  wire _00534_;
  wire _00535_;
  wire _00536_;
  wire _00537_;
  wire _00538_;
  wire _00539_;
  wire _00540_;
  wire _00541_;
  wire _00542_;
  wire _00543_;
  wire _00544_;
  wire _00545_;
  wire _00546_;
  wire _00547_;
  wire _00548_;
  wire _00549_;
  wire _00550_;
  wire _00551_;
  wire _00552_;
  wire _00553_;
  wire _00554_;
  wire _00555_;
  wire _00556_;
  wire _00557_;
  wire _00558_;
  wire _00559_;
  wire _00560_;
  wire _00561_;
  wire _00562_;
  wire _00563_;
  wire _00564_;
  wire _00565_;
  wire _00566_;
  wire _00567_;
  wire _00568_;
  wire _00569_;
  wire _00570_;
  wire _00571_;
  wire _00572_;
  wire _00573_;
  wire _00574_;
  wire _00575_;
  wire _00576_;
  wire _00577_;
  wire _00578_;
  wire _00579_;
  wire _00580_;
  wire _00581_;
  wire _00582_;
  wire _00583_;
  wire _00584_;
  wire _00585_;
  wire _00586_;
  wire _00587_;
  wire _00588_;
  wire _00589_;
  wire _00590_;
  wire _00591_;
  wire _00592_;
  wire _00593_;
  wire _00594_;
  wire _00595_;
  wire _00596_;
  wire _00597_;
  wire _00598_;
  wire _00599_;
  wire _00600_;
  wire _00601_;
  wire _00602_;
  wire _00603_;
  wire _00604_;
  wire _00605_;
  wire _00606_;
  wire _00607_;
  wire _00608_;
  wire _00609_;
  wire _00610_;
  wire _00611_;
  wire _00612_;
  wire _00613_;
  wire _00614_;
  wire _00615_;
  wire _00616_;
  wire _00617_;
  wire _00618_;
  wire _00619_;
  wire _00620_;
  wire _00621_;
  wire _00622_;
  wire _00623_;
  wire _00624_;
  wire _00625_;
  wire _00626_;
  wire _00627_;
  wire _00628_;
  wire _00629_;
  wire _00630_;
  wire _00631_;
  wire _00632_;
  wire _00633_;
  wire _00634_;
  wire _00635_;
  wire _00636_;
  wire _00637_;
  wire _00638_;
  wire _00639_;
  wire _00640_;
  wire _00641_;
  wire _00642_;
  wire _00643_;
  wire _00644_;
  wire _00645_;
  wire _00646_;
  wire _00647_;
  wire _00648_;
  wire _00649_;
  wire _00650_;
  wire _00651_;
  wire _00652_;
  wire _00653_;
  wire _00654_;
  wire _00655_;
  wire _00656_;
  wire _00657_;
  wire _00658_;
  wire _00659_;
  wire _00660_;
  wire _00661_;
  wire _00662_;
  wire _00663_;
  wire _00664_;
  wire _00665_;
  wire _00666_;
  wire _00667_;
  wire _00668_;
  wire _00669_;
  wire _00670_;
  wire _00671_;
  wire _00672_;
  wire _00673_;
  wire _00674_;
  wire _00675_;
  wire _00676_;
  wire _00677_;
  wire _00678_;
  wire _00679_;
  wire _00680_;
  wire _00681_;
  wire _00682_;
  wire _00683_;
  wire _00684_;
  wire _00685_;
  wire _00686_;
  wire _00687_;
  wire _00688_;
  wire _00689_;
  wire _00690_;
  wire _00691_;
  wire _00692_;
  wire _00693_;
  wire _00694_;
  wire _00695_;
  wire _00696_;
  wire _00697_;
  wire _00698_;
  wire _00699_;
  wire _00700_;
  wire _00701_;
  wire _00702_;
  wire _00703_;
  wire _00704_;
  wire _00705_;
  wire _00706_;
  wire _00707_;
  wire _00708_;
  wire _00709_;
  wire _00710_;
  wire _00711_;
  wire _00712_;
  wire _00713_;
  wire _00714_;
  wire _00715_;
  wire _00716_;
  wire _00717_;
  wire _00718_;
  wire _00719_;
  wire _00720_;
  wire _00721_;
  wire _00722_;
  wire _00723_;
  wire _00724_;
  wire _00725_;
  wire _00726_;
  wire _00727_;
  wire _00728_;
  wire _00729_;
  wire _00730_;
  wire _00731_;
  wire _00732_;
  wire _00733_;
  wire _00734_;
  wire _00735_;
  wire _00736_;
  wire _00737_;
  wire _00738_;
  wire _00739_;
  wire _00740_;
  wire _00741_;
  wire _00742_;
  wire _00743_;
  wire _00744_;
  wire _00745_;
  wire _00746_;
  wire _00747_;
  wire _00748_;
  wire _00749_;
  wire _00750_;
  wire _00751_;
  wire _00752_;
  wire _00753_;
  wire _00754_;
  wire _00755_;
  wire _00756_;
  wire _00757_;
  wire _00758_;
  wire _00759_;
  wire _00760_;
  wire _00761_;
  wire _00762_;
  wire _00763_;
  wire _00764_;
  wire _00765_;
  wire _00766_;
  wire _00767_;
  wire _00768_;
  wire _00769_;
  wire _00770_;
  wire _00771_;
  wire _00772_;
  wire _00773_;
  wire _00774_;
  wire _00775_;
  wire _00776_;
  wire _00777_;
  wire _00778_;
  wire _00779_;
  wire _00780_;
  wire _00781_;
  wire _00782_;
  wire _00783_;
  wire _00784_;
  wire _00785_;
  wire _00786_;
  wire _00787_;
  wire _00788_;
  wire _00789_;
  wire _00790_;
  wire _00791_;
  wire _00792_;
  wire _00793_;
  wire _00794_;
  wire _00795_;
  wire _00796_;
  wire _00797_;
  wire _00798_;
  wire _00799_;
  wire _00800_;
  wire _00801_;
  wire _00802_;
  wire _00803_;
  wire _00804_;
  wire _00805_;
  wire _00806_;
  wire _00807_;
  wire _00808_;
  wire _00809_;
  wire _00810_;
  wire _00811_;
  wire _00812_;
  wire _00813_;
  wire _00814_;
  wire _00815_;
  wire _00816_;
  wire _00817_;
  wire _00818_;
  wire _00819_;
  wire _00820_;
  wire _00821_;
  wire _00822_;
  wire _00823_;
  wire _00824_;
  wire _00825_;
  wire _00826_;
  wire _00827_;
  wire _00828_;
  wire _00829_;
  wire _00830_;
  wire _00831_;
  wire _00832_;
  wire _00833_;
  wire _00834_;
  wire _00835_;
  wire _00836_;
  wire _00837_;
  wire _00838_;
  wire _00839_;
  wire _00840_;
  wire _00841_;
  wire _00842_;
  wire _00843_;
  wire _00844_;
  wire _00845_;
  wire _00846_;
  wire _00847_;
  wire _00848_;
  wire _00849_;
  wire _00850_;
  wire _00851_;
  wire _00852_;
  wire _00853_;
  wire _00854_;
  wire _00855_;
  wire _00856_;
  wire _00857_;
  wire _00858_;
  wire _00859_;
  wire _00860_;
  wire _00861_;
  wire _00862_;
  wire _00863_;
  wire _00864_;
  wire _00865_;
  wire _00866_;
  wire _00867_;
  wire _00868_;
  wire _00869_;
  wire _00870_;
  wire _00871_;
  wire _00872_;
  wire _00873_;
  wire _00874_;
  wire _00875_;
  wire _00876_;
  wire _00877_;
  wire _00878_;
  wire _00879_;
  wire _00880_;
  wire _00881_;
  wire _00882_;
  wire _00883_;
  wire _00884_;
  wire _00885_;
  wire _00886_;
  wire _00887_;
  wire _00888_;
  wire _00889_;
  wire _00890_;
  wire _00891_;
  wire _00892_;
  wire _00893_;
  wire _00894_;
  wire _00895_;
  wire _00896_;
  wire _00897_;
  wire _00898_;
  wire _00899_;
  wire _00900_;
  wire _00901_;
  wire _00902_;
  wire _00903_;
  wire _00904_;
  wire _00905_;
  wire _00906_;
  wire _00907_;
  wire _00908_;
  wire _00909_;
  wire _00910_;
  wire _00911_;
  wire _00912_;
  wire _00913_;
  wire _00914_;
  wire _00915_;
  wire _00916_;
  wire _00917_;
  wire _00918_;
  wire _00919_;
  wire _00920_;
  wire _00921_;
  wire _00922_;
  wire _00923_;
  wire _00924_;
  wire _00925_;
  wire _00926_;
  wire _00927_;
  wire _00928_;
  wire _00929_;
  wire _00930_;
  wire _00931_;
  wire _00932_;
  wire _00933_;
  wire _00934_;
  wire _00935_;
  wire _00936_;
  wire _00937_;
  wire _00938_;
  wire _00939_;
  wire _00940_;
  wire _00941_;
  wire _00942_;
  wire _00943_;
  wire _00944_;
  wire _00945_;
  wire _00946_;
  wire _00947_;
  wire _00948_;
  wire _00949_;
  wire _00950_;
  wire _00951_;
  wire _00952_;
  wire _00953_;
  wire _00954_;
  wire _00955_;
  wire _00956_;
  wire _00957_;
  wire _00958_;
  wire _00959_;
  wire _00960_;
  wire _00961_;
  wire _00962_;
  wire _00963_;
  wire _00964_;
  wire _00965_;
  wire _00966_;
  wire _00967_;
  wire _00968_;
  wire _00969_;
  wire _00970_;
  wire _00971_;
  wire _00972_;
  wire _00973_;
  wire _00974_;
  wire _00975_;
  wire _00976_;
  wire _00977_;
  wire _00978_;
  wire _00979_;
  wire _00980_;
  wire _00981_;
  wire _00982_;
  wire _00983_;
  wire _00984_;
  wire _00985_;
  wire _00986_;
  wire _00987_;
  wire _00988_;
  wire _00989_;
  wire _00990_;
  wire _00991_;
  wire _00992_;
  wire _00993_;
  wire _00994_;
  wire _00995_;
  wire _00996_;
  wire _00997_;
  wire _00998_;
  wire _00999_;
  wire _01000_;
  wire _01001_;
  wire _01002_;
  wire _01003_;
  wire _01004_;
  wire _01005_;
  wire _01006_;
  wire _01007_;
  wire _01008_;
  wire _01009_;
  wire _01010_;
  wire _01011_;
  wire _01012_;
  wire _01013_;
  wire _01014_;
  wire _01015_;
  wire _01016_;
  wire _01017_;
  wire _01018_;
  wire _01019_;
  wire _01020_;
  wire _01021_;
  wire _01022_;
  wire _01023_;
  wire _01024_;
  wire _01025_;
  wire _01026_;
  wire _01027_;
  wire _01028_;
  wire _01029_;
  wire _01030_;
  wire _01031_;
  wire _01032_;
  wire _01033_;
  wire _01034_;
  wire _01035_;
  wire _01036_;
  wire _01037_;
  wire _01038_;
  wire _01039_;
  wire _01040_;
  wire _01041_;
  wire _01042_;
  wire _01043_;
  wire _01044_;
  wire _01045_;
  wire _01046_;
  wire _01047_;
  wire _01048_;
  wire _01049_;
  wire _01050_;
  wire _01051_;
  wire _01052_;
  wire _01053_;
  wire _01054_;
  wire _01055_;
  wire _01056_;
  wire _01057_;
  wire _01058_;
  wire _01059_;
  wire _01060_;
  wire _01061_;
  wire _01062_;
  wire _01063_;
  wire _01064_;
  wire _01065_;
  wire _01066_;
  wire _01067_;
  wire _01068_;
  wire _01069_;
  wire _01070_;
  wire _01071_;
  wire _01072_;
  wire _01073_;
  wire _01074_;
  wire _01075_;
  wire _01076_;
  wire _01077_;
  wire _01078_;
  wire _01079_;
  wire _01080_;
  wire _01081_;
  wire _01082_;
  wire _01083_;
  wire _01084_;
  wire _01085_;
  wire _01086_;
  wire _01087_;
  wire _01088_;
  wire _01089_;
  wire _01090_;
  wire _01091_;
  wire _01092_;
  wire _01093_;
  wire _01094_;
  wire _01095_;
  wire _01096_;
  wire _01097_;
  wire _01098_;
  wire _01099_;
  wire _01100_;
  wire _01101_;
  wire _01102_;
  wire _01103_;
  wire _01104_;
  wire _01105_;
  wire _01106_;
  wire _01107_;
  wire _01108_;
  wire _01109_;
  wire _01110_;
  wire _01111_;
  wire _01112_;
  wire _01113_;
  wire _01114_;
  wire _01115_;
  wire _01116_;
  wire _01117_;
  wire _01118_;
  wire _01119_;
  wire _01120_;
  wire _01121_;
  wire _01122_;
  wire _01123_;
  wire _01124_;
  wire _01125_;
  wire _01126_;
  wire _01127_;
  wire _01128_;
  wire _01129_;
  wire _01130_;
  wire _01131_;
  wire _01132_;
  wire _01133_;
  wire _01134_;
  wire _01135_;
  wire _01136_;
  wire _01137_;
  wire _01138_;
  wire _01139_;
  wire _01140_;
  wire _01141_;
  wire _01142_;
  wire _01143_;
  wire _01144_;
  wire _01145_;
  wire _01146_;
  wire _01147_;
  wire _01148_;
  wire _01149_;
  wire _01150_;
  wire _01151_;
  wire _01152_;
  wire _01153_;
  wire _01154_;
  wire _01155_;
  wire _01156_;
  wire _01157_;
  wire _01158_;
  wire _01159_;
  wire _01160_;
  wire _01161_;
  wire _01162_;
  wire _01163_;
  wire _01164_;
  wire _01165_;
  wire _01166_;
  wire _01167_;
  wire _01168_;
  wire _01169_;
  wire _01170_;
  wire _01171_;
  wire _01172_;
  wire _01173_;
  wire _01174_;
  wire _01175_;
  wire _01176_;
  wire _01177_;
  wire _01178_;
  wire _01179_;
  wire _01180_;
  wire _01181_;
  wire _01182_;
  wire _01183_;
  wire _01184_;
  wire _01185_;
  wire _01186_;
  wire _01187_;
  wire _01188_;
  wire _01189_;
  wire _01190_;
  wire _01191_;
  wire _01192_;
  wire _01193_;
  wire _01194_;
  wire _01195_;
  wire _01196_;
  wire _01197_;
  wire _01198_;
  wire _01199_;
  wire _01200_;
  wire _01201_;
  wire _01202_;
  wire _01203_;
  wire _01204_;
  wire _01205_;
  wire _01206_;
  wire _01207_;
  wire _01208_;
  wire _01209_;
  wire _01210_;
  wire _01211_;
  wire _01212_;
  wire _01213_;
  wire _01214_;
  wire _01215_;
  wire _01216_;
  wire _01217_;
  wire _01218_;
  wire _01219_;
  wire _01220_;
  wire _01221_;
  wire _01222_;
  wire _01223_;
  wire _01224_;
  wire _01225_;
  wire _01226_;
  wire _01227_;
  wire _01228_;
  wire _01229_;
  wire _01230_;
  wire _01231_;
  wire _01232_;
  wire _01233_;
  wire _01234_;
  wire _01235_;
  wire _01236_;
  wire _01237_;
  wire _01238_;
  wire _01239_;
  wire _01240_;
  wire _01241_;
  wire _01242_;
  wire _01243_;
  wire _01244_;
  wire _01245_;
  wire _01246_;
  wire _01247_;
  wire _01248_;
  wire _01249_;
  wire _01250_;
  wire _01251_;
  wire _01252_;
  wire _01253_;
  wire _01254_;
  wire _01255_;
  wire _01256_;
  wire _01257_;
  wire _01258_;
  wire _01259_;
  wire _01260_;
  wire _01261_;
  wire _01262_;
  wire _01263_;
  wire _01264_;
  wire _01265_;
  wire _01266_;
  wire _01267_;
  wire _01268_;
  wire _01269_;
  wire _01270_;
  wire _01271_;
  wire _01272_;
  wire _01273_;
  wire _01274_;
  wire _01275_;
  wire _01276_;
  wire _01277_;
  wire _01278_;
  wire _01279_;
  wire _01280_;
  wire _01281_;
  wire _01282_;
  wire _01283_;
  wire _01284_;
  wire _01285_;
  wire _01286_;
  wire _01287_;
  wire _01288_;
  wire _01289_;
  wire _01290_;
  wire _01291_;
  wire _01292_;
  wire _01293_;
  wire _01294_;
  wire _01295_;
  wire _01296_;
  wire _01297_;
  wire _01298_;
  wire _01299_;
  wire _01300_;
  wire _01301_;
  wire _01302_;
  wire _01303_;
  wire _01304_;
  wire _01305_;
  wire _01306_;
  wire _01307_;
  wire _01308_;
  wire _01309_;
  wire _01310_;
  wire _01311_;
  wire _01312_;
  wire _01313_;
  wire _01314_;
  wire _01315_;
  wire _01316_;
  wire _01317_;
  wire _01318_;
  wire _01319_;
  wire _01320_;
  wire _01321_;
  wire _01322_;
  wire _01323_;
  wire _01324_;
  wire _01325_;
  wire _01326_;
  wire _01327_;
  wire _01328_;
  wire _01329_;
  wire _01330_;
  wire _01331_;
  wire _01332_;
  wire _01333_;
  wire _01334_;
  wire _01335_;
  wire _01336_;
  wire _01337_;
  wire _01338_;
  wire _01339_;
  wire _01340_;
  wire _01341_;
  wire _01342_;
  wire _01343_;
  wire _01344_;
  wire _01345_;
  wire _01346_;
  wire _01347_;
  wire _01348_;
  wire _01349_;
  wire _01350_;
  wire _01351_;
  wire _01352_;
  wire _01353_;
  wire _01354_;
  wire _01355_;
  wire _01356_;
  wire _01357_;
  wire _01358_;
  wire _01359_;
  wire _01360_;
  wire _01361_;
  wire _01362_;
  wire _01363_;
  wire _01364_;
  wire _01365_;
  wire _01366_;
  wire _01367_;
  wire _01368_;
  wire _01369_;
  wire _01370_;
  wire _01371_;
  wire _01372_;
  wire _01373_;
  wire _01374_;
  wire _01375_;
  wire _01376_;
  wire _01377_;
  wire _01378_;
  wire _01379_;
  wire _01380_;
  wire _01381_;
  wire _01382_;
  wire _01383_;
  wire _01384_;
  wire _01385_;
  wire _01386_;
  wire _01387_;
  wire _01388_;
  wire _01389_;
  wire _01390_;
  wire _01391_;
  wire _01392_;
  wire _01393_;
  wire _01394_;
  wire _01395_;
  wire _01396_;
  wire _01397_;
  wire _01398_;
  wire _01399_;
  wire _01400_;
  wire _01401_;
  wire _01402_;
  wire _01403_;
  wire _01404_;
  wire _01405_;
  wire _01406_;
  wire _01407_;
  wire _01408_;
  wire _01409_;
  wire _01410_;
  wire _01411_;
  wire _01412_;
  wire _01413_;
  wire _01414_;
  wire _01415_;
  wire _01416_;
  wire _01417_;
  wire _01418_;
  wire _01419_;
  wire _01420_;
  wire _01421_;
  wire _01422_;
  wire _01423_;
  wire _01424_;
  wire _01425_;
  wire _01426_;
  wire _01427_;
  wire _01428_;
  wire _01429_;
  wire _01430_;
  wire _01431_;
  wire _01432_;
  wire _01433_;
  wire _01434_;
  wire _01435_;
  wire _01436_;
  wire _01437_;
  wire _01438_;
  wire _01439_;
  wire _01440_;
  wire _01441_;
  wire _01442_;
  wire _01443_;
  wire _01444_;
  wire _01445_;
  wire _01446_;
  wire _01447_;
  wire _01448_;
  wire _01449_;
  wire _01450_;
  wire _01451_;
  wire _01452_;
  wire _01453_;
  wire _01454_;
  wire _01455_;
  wire _01456_;
  wire _01457_;
  wire _01458_;
  wire _01459_;
  wire _01460_;
  wire _01461_;
  wire _01462_;
  wire _01463_;
  wire _01464_;
  wire _01465_;
  wire _01466_;
  wire _01467_;
  wire _01468_;
  wire _01469_;
  wire _01470_;
  wire _01471_;
  wire _01472_;
  wire _01473_;
  wire _01474_;
  wire _01475_;
  wire _01476_;
  wire _01477_;
  wire _01478_;
  wire _01479_;
  wire _01480_;
  wire _01481_;
  wire _01482_;
  wire _01483_;
  wire _01484_;
  wire _01485_;
  wire _01486_;
  wire _01487_;
  wire _01488_;
  wire _01489_;
  wire _01490_;
  wire _01491_;
  wire _01492_;
  wire _01493_;
  wire _01494_;
  wire _01495_;
  wire _01496_;
  wire _01497_;
  wire _01498_;
  wire _01499_;
  wire _01500_;
  wire _01501_;
  wire _01502_;
  wire _01503_;
  wire _01504_;
  wire _01505_;
  wire _01506_;
  wire _01507_;
  wire _01508_;
  wire _01509_;
  wire _01510_;
  wire _01511_;
  wire _01512_;
  wire _01513_;
  wire _01514_;
  wire _01515_;
  wire _01516_;
  wire _01517_;
  wire _01518_;
  wire _01519_;
  wire _01520_;
  wire _01521_;
  wire _01522_;
  wire _01523_;
  wire _01524_;
  wire _01525_;
  wire _01526_;
  wire _01527_;
  wire _01528_;
  wire _01529_;
  wire _01530_;
  wire _01531_;
  wire _01532_;
  wire _01533_;
  wire _01534_;
  wire _01535_;
  wire _01536_;
  wire _01537_;
  wire _01538_;
  wire _01539_;
  wire _01540_;
  wire _01541_;
  wire _01542_;
  wire _01543_;
  wire _01544_;
  wire _01545_;
  wire _01546_;
  wire _01547_;
  wire _01548_;
  wire _01549_;
  wire _01550_;
  wire _01551_;
  wire _01552_;
  wire _01553_;
  wire _01554_;
  wire _01555_;
  wire _01556_;
  wire _01557_;
  wire _01558_;
  wire _01559_;
  wire _01560_;
  wire _01561_;
  wire _01562_;
  wire _01563_;
  wire _01564_;
  wire _01565_;
  wire _01566_;
  wire _01567_;
  wire _01568_;
  wire _01569_;
  wire _01570_;
  wire _01571_;
  wire _01572_;
  wire _01573_;
  wire _01574_;
  wire _01575_;
  wire _01576_;
  wire _01577_;
  wire _01578_;
  wire _01579_;
  wire _01580_;
  wire _01581_;
  wire _01582_;
  wire _01583_;
  wire _01584_;
  wire _01585_;
  wire _01586_;
  wire _01587_;
  wire _01588_;
  wire _01589_;
  wire _01590_;
  wire _01591_;
  wire _01592_;
  wire _01593_;
  wire _01594_;
  wire _01595_;
  wire _01596_;
  wire _01597_;
  wire _01598_;
  wire _01599_;
  wire _01600_;
  wire _01601_;
  wire _01602_;
  wire _01603_;
  wire _01604_;
  wire _01605_;
  wire _01606_;
  wire _01607_;
  wire _01608_;
  wire _01609_;
  wire _01610_;
  wire _01611_;
  wire _01612_;
  wire _01613_;
  wire _01614_;
  wire _01615_;
  wire _01616_;
  wire _01617_;
  wire _01618_;
  wire _01619_;
  wire _01620_;
  wire _01621_;
  wire _01622_;
  wire _01623_;
  wire _01624_;
  wire _01625_;
  wire _01626_;
  wire _01627_;
  wire _01628_;
  wire _01629_;
  wire _01630_;
  wire _01631_;
  wire _01632_;
  wire _01633_;
  wire _01634_;
  wire _01635_;
  wire _01636_;
  wire _01637_;
  wire _01638_;
  wire _01639_;
  wire _01640_;
  wire _01641_;
  wire _01642_;
  wire _01643_;
  wire _01644_;
  wire _01645_;
  wire _01646_;
  wire _01647_;
  wire _01648_;
  wire _01649_;
  wire _01650_;
  wire _01651_;
  wire _01652_;
  wire _01653_;
  wire _01654_;
  wire _01655_;
  wire _01656_;
  wire _01657_;
  wire _01658_;
  wire _01659_;
  wire _01660_;
  wire _01661_;
  wire _01662_;
  wire _01663_;
  wire _01664_;
  wire _01665_;
  wire _01666_;
  wire _01667_;
  wire _01668_;
  wire _01669_;
  wire _01670_;
  wire _01671_;
  wire _01672_;
  wire _01673_;
  wire _01674_;
  wire _01675_;
  wire _01676_;
  wire _01677_;
  wire _01678_;
  wire _01679_;
  wire _01680_;
  wire _01681_;
  wire _01682_;
  wire _01683_;
  wire _01684_;
  wire _01685_;
  wire _01686_;
  wire _01687_;
  wire _01688_;
  wire _01689_;
  wire _01690_;
  wire _01691_;
  wire _01692_;
  wire _01693_;
  wire _01694_;
  wire _01695_;
  wire _01696_;
  wire _01697_;
  wire _01698_;
  wire _01699_;
  wire _01700_;
  wire _01701_;
  wire _01702_;
  wire _01703_;
  wire _01704_;
  wire _01705_;
  wire _01706_;
  wire _01707_;
  wire _01708_;
  wire _01709_;
  wire _01710_;
  wire _01711_;
  wire _01712_;
  wire _01713_;
  wire _01714_;
  wire _01715_;
  wire _01716_;
  wire _01717_;
  wire _01718_;
  wire _01719_;
  wire _01720_;
  wire _01721_;
  wire _01722_;
  wire _01723_;
  wire _01724_;
  wire _01725_;
  wire _01726_;
  wire _01727_;
  wire _01728_;
  wire _01729_;
  wire _01730_;
  wire _01731_;
  wire _01732_;
  wire _01733_;
  wire _01734_;
  wire _01735_;
  wire _01736_;
  wire _01737_;
  wire _01738_;
  wire _01739_;
  wire _01740_;
  wire _01741_;
  wire _01742_;
  wire _01743_;
  wire _01744_;
  wire _01745_;
  wire _01746_;
  wire _01747_;
  wire _01748_;
  wire _01749_;
  wire _01750_;
  wire _01751_;
  wire _01752_;
  wire _01753_;
  wire _01754_;
  wire _01755_;
  wire _01756_;
  wire _01757_;
  wire _01758_;
  wire _01759_;
  wire _01760_;
  wire _01761_;
  wire _01762_;
  wire _01763_;
  wire _01764_;
  wire _01765_;
  wire _01766_;
  wire _01767_;
  wire _01768_;
  wire _01769_;
  wire _01770_;
  wire _01771_;
  wire _01772_;
  wire _01773_;
  wire _01774_;
  wire _01775_;
  wire _01776_;
  wire _01777_;
  wire _01778_;
  wire _01779_;
  wire _01780_;
  wire _01781_;
  wire _01782_;
  wire _01783_;
  wire _01784_;
  wire _01785_;
  wire _01786_;
  wire _01787_;
  wire _01788_;
  wire _01789_;
  wire _01790_;
  wire _01791_;
  wire _01792_;
  wire _01793_;
  wire _01794_;
  wire _01795_;
  wire _01796_;
  wire _01797_;
  wire _01798_;
  wire _01799_;
  wire _01800_;
  wire _01801_;
  wire _01802_;
  wire _01803_;
  wire _01804_;
  wire _01805_;
  wire _01806_;
  wire _01807_;
  wire _01808_;
  wire _01809_;
  wire _01810_;
  wire _01811_;
  wire _01812_;
  wire _01813_;
  wire _01814_;
  wire _01815_;
  wire _01816_;
  wire _01817_;
  wire _01818_;
  wire _01819_;
  wire _01820_;
  wire _01821_;
  wire _01822_;
  wire _01823_;
  wire _01824_;
  wire _01825_;
  wire _01826_;
  wire _01827_;
  wire _01828_;
  wire _01829_;
  wire _01830_;
  wire _01831_;
  wire _01832_;
  wire _01833_;
  wire _01834_;
  wire _01835_;
  wire _01836_;
  wire _01837_;
  wire _01838_;
  wire _01839_;
  wire _01840_;
  wire _01841_;
  wire _01842_;
  wire _01843_;
  wire _01844_;
  wire _01845_;
  wire _01846_;
  wire _01847_;
  wire _01848_;
  wire _01849_;
  wire _01850_;
  wire _01851_;
  wire _01852_;
  wire _01853_;
  wire _01854_;
  wire _01855_;
  wire _01856_;
  wire _01857_;
  wire _01858_;
  wire _01859_;
  wire _01860_;
  wire _01861_;
  wire _01862_;
  wire _01863_;
  wire _01864_;
  wire _01865_;
  wire _01866_;
  wire _01867_;
  wire _01868_;
  wire _01869_;
  wire _01870_;
  wire _01871_;
  wire _01872_;
  wire _01873_;
  wire _01874_;
  wire _01875_;
  wire _01876_;
  wire _01877_;
  wire _01878_;
  wire _01879_;
  wire _01880_;
  wire _01881_;
  wire _01882_;
  wire _01883_;
  wire _01884_;
  wire _01885_;
  wire _01886_;
  wire _01887_;
  wire _01888_;
  wire _01889_;
  wire _01890_;
  wire _01891_;
  wire _01892_;
  wire _01893_;
  wire _01894_;
  wire _01895_;
  wire _01896_;
  wire _01897_;
  wire _01898_;
  wire _01899_;
  wire _01900_;
  wire _01901_;
  wire _01902_;
  wire _01903_;
  wire _01904_;
  wire _01905_;
  wire _01906_;
  wire _01907_;
  wire _01908_;
  wire _01909_;
  wire _01910_;
  wire _01911_;
  wire _01912_;
  wire _01913_;
  wire _01914_;
  wire _01915_;
  wire _01916_;
  wire _01917_;
  wire _01918_;
  wire _01919_;
  wire _01920_;
  wire _01921_;
  wire _01922_;
  wire _01923_;
  wire _01924_;
  wire _01925_;
  wire _01926_;
  wire _01927_;
  wire _01928_;
  wire _01929_;
  wire _01930_;
  wire _01931_;
  wire _01932_;
  wire _01933_;
  wire _01934_;
  wire _01935_;
  wire _01936_;
  wire _01937_;
  wire _01938_;
  wire _01939_;
  wire _01940_;
  wire _01941_;
  wire _01942_;
  wire _01943_;
  wire _01944_;
  wire _01945_;
  wire _01946_;
  wire _01947_;
  wire _01948_;
  wire _01949_;
  wire _01950_;
  wire _01951_;
  wire _01952_;
  wire _01953_;
  wire _01954_;
  wire _01955_;
  wire _01956_;
  wire _01957_;
  wire _01958_;
  wire _01959_;
  wire _01960_;
  wire _01961_;
  wire _01962_;
  wire _01963_;
  wire _01964_;
  wire _01965_;
  wire _01966_;
  wire _01967_;
  wire _01968_;
  wire _01969_;
  wire _01970_;
  wire _01971_;
  wire _01972_;
  wire _01973_;
  wire _01974_;
  wire _01975_;
  wire _01976_;
  wire _01977_;
  wire _01978_;
  wire _01979_;
  wire _01980_;
  wire _01981_;
  wire _01982_;
  wire _01983_;
  wire _01984_;
  wire _01985_;
  wire _01986_;
  wire _01987_;
  wire _01988_;
  wire _01989_;
  wire _01990_;
  wire _01991_;
  wire _01992_;
  wire _01993_;
  wire _01994_;
  wire _01995_;
  wire _01996_;
  wire _01997_;
  wire _01998_;
  wire _01999_;
  wire _02000_;
  wire _02001_;
  wire _02002_;
  wire _02003_;
  wire _02004_;
  wire _02005_;
  wire _02006_;
  wire _02007_;
  wire _02008_;
  wire _02009_;
  wire _02010_;
  wire _02011_;
  wire _02012_;
  wire _02013_;
  wire _02014_;
  wire _02015_;
  wire _02016_;
  wire _02017_;
  wire _02018_;
  wire _02019_;
  wire _02020_;
  wire _02021_;
  wire _02022_;
  wire _02023_;
  wire _02024_;
  wire _02025_;
  wire _02026_;
  wire _02027_;
  wire _02028_;
  wire _02029_;
  wire _02030_;
  wire _02031_;
  wire _02032_;
  wire _02033_;
  wire _02034_;
  wire _02035_;
  wire _02036_;
  wire _02037_;
  wire _02038_;
  wire _02039_;
  wire _02040_;
  wire _02041_;
  wire _02042_;
  wire _02043_;
  wire _02044_;
  wire _02045_;
  wire _02046_;
  wire _02047_;
  wire _02048_;
  wire _02049_;
  wire _02050_;
  wire _02051_;
  wire _02052_;
  wire _02053_;
  wire _02054_;
  wire _02055_;
  wire _02056_;
  wire _02057_;
  wire _02058_;
  wire _02059_;
  wire _02060_;
  wire _02061_;
  wire _02062_;
  wire _02063_;
  wire _02064_;
  wire _02065_;
  wire _02066_;
  wire _02067_;
  wire _02068_;
  wire _02069_;
  wire _02070_;
  wire _02071_;
  wire _02072_;
  wire _02073_;
  wire _02074_;
  wire _02075_;
  wire _02076_;
  wire _02077_;
  wire _02078_;
  wire _02079_;
  wire _02080_;
  wire _02081_;
  wire _02082_;
  wire _02083_;
  wire _02084_;
  wire _02085_;
  wire _02086_;
  wire _02087_;
  wire _02088_;
  wire _02089_;
  wire _02090_;
  wire _02091_;
  wire _02092_;
  wire _02093_;
  wire _02094_;
  wire _02095_;
  wire _02096_;
  wire _02097_;
  wire _02098_;
  wire _02099_;
  wire _02100_;
  wire _02101_;
  wire _02102_;
  wire _02103_;
  wire _02104_;
  wire _02105_;
  wire _02106_;
  wire _02107_;
  wire _02108_;
  wire _02109_;
  wire _02110_;
  wire _02111_;
  wire _02112_;
  wire _02113_;
  wire _02114_;
  wire _02115_;
  wire _02116_;
  wire _02117_;
  wire _02118_;
  wire _02119_;
  wire _02120_;
  wire _02121_;
  wire _02122_;
  wire _02123_;
  wire _02124_;
  wire _02125_;
  wire _02126_;
  wire _02127_;
  wire _02128_;
  wire _02129_;
  wire _02130_;
  wire _02131_;
  wire _02132_;
  wire _02133_;
  wire _02134_;
  wire _02135_;
  wire _02136_;
  wire _02137_;
  wire _02138_;
  wire _02139_;
  wire _02140_;
  wire _02141_;
  wire _02142_;
  wire _02143_;
  wire _02144_;
  wire _02145_;
  wire _02146_;
  wire _02147_;
  wire _02148_;
  wire _02149_;
  wire _02150_;
  wire _02151_;
  wire _02152_;
  wire _02153_;
  wire _02154_;
  wire _02155_;
  wire _02156_;
  wire _02157_;
  wire _02158_;
  wire _02159_;
  wire _02160_;
  wire _02161_;
  wire _02162_;
  wire _02163_;
  wire _02164_;
  wire _02165_;
  wire _02166_;
  wire _02167_;
  wire _02168_;
  wire _02169_;
  wire _02170_;
  wire _02171_;
  wire _02172_;
  wire _02173_;
  wire _02174_;
  wire _02175_;
  wire _02176_;
  wire _02177_;
  wire _02178_;
  wire _02179_;
  wire _02180_;
  wire _02181_;
  wire _02182_;
  wire _02183_;
  wire _02184_;
  wire _02185_;
  wire _02186_;
  wire _02187_;
  wire _02188_;
  wire _02189_;
  wire _02190_;
  wire _02191_;
  wire _02192_;
  wire _02193_;
  wire _02194_;
  wire _02195_;
  wire _02196_;
  wire _02197_;
  wire _02198_;
  wire _02199_;
  wire _02200_;
  wire _02201_;
  wire _02202_;
  wire _02203_;
  wire _02204_;
  wire _02205_;
  wire _02206_;
  wire _02207_;
  wire _02208_;
  wire _02209_;
  wire _02210_;
  wire _02211_;
  wire _02212_;
  wire _02213_;
  wire _02214_;
  wire _02215_;
  wire _02216_;
  wire _02217_;
  wire _02218_;
  wire _02219_;
  wire _02220_;
  wire _02221_;
  wire _02222_;
  wire _02223_;
  wire _02224_;
  wire _02225_;
  wire _02226_;
  wire _02227_;
  wire _02228_;
  wire _02229_;
  wire _02230_;
  wire _02231_;
  wire _02232_;
  wire _02233_;
  wire _02234_;
  wire _02235_;
  wire _02236_;
  wire _02237_;
  wire _02238_;
  wire _02239_;
  wire _02240_;
  wire _02241_;
  wire _02242_;
  wire _02243_;
  wire _02244_;
  wire _02245_;
  wire _02246_;
  wire _02247_;
  wire _02248_;
  wire _02249_;
  wire _02250_;
  wire _02251_;
  wire _02252_;
  wire _02253_;
  wire _02254_;
  wire _02255_;
  wire _02256_;
  wire _02257_;
  wire _02258_;
  wire _02259_;
  wire _02260_;
  wire _02261_;
  wire _02262_;
  wire _02263_;
  wire _02264_;
  wire _02265_;
  wire _02266_;
  wire _02267_;
  wire _02268_;
  wire _02269_;
  wire _02270_;
  wire _02271_;
  wire _02272_;
  wire _02273_;
  wire _02274_;
  wire _02275_;
  wire _02276_;
  wire _02277_;
  wire _02278_;
  wire _02279_;
  wire _02280_;
  wire _02281_;
  wire _02282_;
  wire _02283_;
  wire _02284_;
  wire _02285_;
  wire _02286_;
  wire _02287_;
  wire _02288_;
  wire _02289_;
  wire _02290_;
  wire _02291_;
  wire _02292_;
  wire _02293_;
  wire _02294_;
  wire _02295_;
  wire _02296_;
  wire _02297_;
  wire _02298_;
  wire _02299_;
  wire _02300_;
  wire _02301_;
  wire _02302_;
  wire _02303_;
  wire _02304_;
  wire _02305_;
  wire _02306_;
  wire _02307_;
  wire _02308_;
  wire _02309_;
  wire _02310_;
  wire _02311_;
  wire _02312_;
  wire _02313_;
  wire _02314_;
  wire _02315_;
  wire _02316_;
  wire _02317_;
  wire _02318_;
  wire _02319_;
  wire _02320_;
  wire _02321_;
  wire _02322_;
  wire _02323_;
  wire _02324_;
  wire _02325_;
  wire _02326_;
  wire _02327_;
  wire _02328_;
  wire _02329_;
  wire _02330_;
  wire _02331_;
  wire _02332_;
  wire _02333_;
  wire _02334_;
  wire _02335_;
  wire _02336_;
  wire _02337_;
  wire _02338_;
  wire _02339_;
  wire _02340_;
  wire _02341_;
  wire _02342_;
  wire _02343_;
  wire _02344_;
  wire _02345_;
  wire _02346_;
  wire _02347_;
  wire _02348_;
  wire _02349_;
  wire _02350_;
  wire _02351_;
  wire _02352_;
  wire _02353_;
  wire _02354_;
  wire _02355_;
  wire _02356_;
  wire _02357_;
  wire _02358_;
  wire _02359_;
  wire _02360_;
  wire _02361_;
  wire _02362_;
  wire _02363_;
  wire _02364_;
  wire _02365_;
  wire _02366_;
  wire _02367_;
  wire _02368_;
  wire _02369_;
  wire _02370_;
  wire _02371_;
  wire _02372_;
  wire _02373_;
  wire _02374_;
  wire _02375_;
  wire _02376_;
  wire _02377_;
  wire _02378_;
  wire _02379_;
  wire _02380_;
  wire _02381_;
  wire _02382_;
  wire _02383_;
  wire _02384_;
  wire _02385_;
  wire _02386_;
  wire _02387_;
  wire _02388_;
  wire _02389_;
  wire _02390_;
  wire _02391_;
  wire _02392_;
  wire _02393_;
  wire _02394_;
  wire _02395_;
  wire _02396_;
  wire _02397_;
  wire _02398_;
  wire _02399_;
  wire _02400_;
  wire _02401_;
  wire _02402_;
  wire _02403_;
  wire _02404_;
  wire _02405_;
  wire _02406_;
  wire _02407_;
  wire _02408_;
  wire _02409_;
  wire _02410_;
  wire _02411_;
  wire _02412_;
  wire _02413_;
  wire _02414_;
  wire _02415_;
  wire _02416_;
  wire _02417_;
  wire _02418_;
  wire _02419_;
  wire _02420_;
  wire _02421_;
  wire _02422_;
  wire _02423_;
  wire _02424_;
  wire _02425_;
  wire _02426_;
  wire _02427_;
  wire _02428_;
  wire _02429_;
  wire _02430_;
  wire _02431_;
  wire _02432_;
  wire _02433_;
  wire _02434_;
  wire _02435_;
  wire _02436_;
  wire _02437_;
  wire _02438_;
  wire _02439_;
  wire _02440_;
  wire _02441_;
  wire _02442_;
  wire _02443_;
  wire _02444_;
  wire _02445_;
  wire _02446_;
  wire _02447_;
  wire _02448_;
  wire _02449_;
  wire _02450_;
  wire _02451_;
  wire _02452_;
  wire _02453_;
  wire _02454_;
  wire _02455_;
  wire _02456_;
  wire _02457_;
  wire _02458_;
  wire _02459_;
  wire _02460_;
  wire _02461_;
  wire _02462_;
  wire _02463_;
  wire _02464_;
  wire _02465_;
  wire _02466_;
  wire _02467_;
  wire _02468_;
  wire _02469_;
  wire _02470_;
  wire _02471_;
  wire _02472_;
  wire _02473_;
  wire _02474_;
  wire _02475_;
  wire _02476_;
  wire _02477_;
  wire _02478_;
  wire _02479_;
  wire _02480_;
  wire _02481_;
  wire _02482_;
  wire _02483_;
  wire _02484_;
  wire _02485_;
  wire _02486_;
  wire _02487_;
  wire _02488_;
  wire _02489_;
  wire _02490_;
  wire _02491_;
  wire _02492_;
  wire _02493_;
  wire _02494_;
  wire _02495_;
  wire _02496_;
  wire _02497_;
  wire _02498_;
  wire _02499_;
  wire _02500_;
  wire _02501_;
  wire _02502_;
  wire _02503_;
  wire _02504_;
  wire _02505_;
  wire _02506_;
  wire _02507_;
  wire _02508_;
  wire _02509_;
  wire _02510_;
  wire _02511_;
  wire _02512_;
  wire _02513_;
  wire _02514_;
  wire _02515_;
  wire _02516_;
  wire _02517_;
  wire _02518_;
  wire _02519_;
  wire _02520_;
  wire _02521_;
  wire _02522_;
  wire _02523_;
  wire _02524_;
  wire _02525_;
  wire _02526_;
  wire _02527_;
  wire _02528_;
  wire _02529_;
  wire _02530_;
  wire _02531_;
  wire _02532_;
  wire _02533_;
  wire _02534_;
  wire _02535_;
  wire _02536_;
  wire _02537_;
  wire _02538_;
  wire _02539_;
  wire _02540_;
  wire _02541_;
  wire _02542_;
  wire _02543_;
  wire _02544_;
  wire _02545_;
  wire _02546_;
  wire _02547_;
  wire _02548_;
  wire _02549_;
  wire _02550_;
  wire _02551_;
  wire _02552_;
  wire _02553_;
  wire _02554_;
  wire _02555_;
  wire _02556_;
  wire _02557_;
  wire _02558_;
  wire _02559_;
  wire _02560_;
  wire _02561_;
  wire _02562_;
  wire _02563_;
  wire _02564_;
  wire _02565_;
  wire _02566_;
  wire _02567_;
  wire _02568_;
  wire _02569_;
  wire _02570_;
  wire _02571_;
  wire _02572_;
  wire _02573_;
  wire _02574_;
  wire _02575_;
  wire _02576_;
  wire _02577_;
  wire _02578_;
  wire _02579_;
  wire _02580_;
  wire _02581_;
  wire _02582_;
  wire _02583_;
  wire _02584_;
  wire _02585_;
  wire _02586_;
  wire _02587_;
  wire _02588_;
  wire _02589_;
  wire _02590_;
  wire _02591_;
  wire _02592_;
  wire _02593_;
  wire _02594_;
  wire _02595_;
  wire _02596_;
  wire _02597_;
  wire _02598_;
  wire _02599_;
  wire _02600_;
  wire _02601_;
  wire _02602_;
  wire _02603_;
  wire _02604_;
  wire _02605_;
  wire _02606_;
  wire _02607_;
  wire _02608_;
  wire _02609_;
  wire _02610_;
  wire _02611_;
  wire _02612_;
  wire _02613_;
  wire _02614_;
  wire _02615_;
  wire _02616_;
  wire _02617_;
  wire _02618_;
  wire _02619_;
  wire _02620_;
  wire _02621_;
  wire _02622_;
  wire _02623_;
  wire _02624_;
  wire _02625_;
  wire _02626_;
  wire _02627_;
  wire _02628_;
  wire _02629_;
  wire _02630_;
  wire _02631_;
  wire _02632_;
  wire _02633_;
  wire _02634_;
  wire _02635_;
  wire _02636_;
  wire _02637_;
  wire _02638_;
  wire _02639_;
  wire _02640_;
  wire _02641_;
  wire _02642_;
  wire _02643_;
  wire _02644_;
  wire _02645_;
  wire _02646_;
  wire _02647_;
  wire _02648_;
  wire _02649_;
  wire _02650_;
  wire _02651_;
  wire _02652_;
  wire _02653_;
  wire _02654_;
  wire _02655_;
  wire _02656_;
  wire _02657_;
  wire _02658_;
  wire _02659_;
  wire _02660_;
  wire _02661_;
  wire _02662_;
  wire _02663_;
  wire _02664_;
  wire _02665_;
  wire _02666_;
  wire _02667_;
  wire _02668_;
  wire _02669_;
  wire _02670_;
  wire _02671_;
  wire _02672_;
  wire _02673_;
  wire _02674_;
  wire _02675_;
  wire _02676_;
  wire _02677_;
  wire _02678_;
  wire _02679_;
  wire _02680_;
  wire _02681_;
  wire _02682_;
  wire _02683_;
  wire _02684_;
  wire _02685_;
  wire _02686_;
  wire _02687_;
  wire _02688_;
  wire _02689_;
  wire _02690_;
  wire _02691_;
  wire _02692_;
  wire _02693_;
  wire _02694_;
  wire _02695_;
  wire _02696_;
  wire _02697_;
  wire _02698_;
  wire _02699_;
  wire _02700_;
  wire _02701_;
  wire _02702_;
  wire _02703_;
  wire _02704_;
  wire _02705_;
  wire _02706_;
  wire _02707_;
  wire _02708_;
  wire _02709_;
  wire _02710_;
  wire _02711_;
  wire _02712_;
  wire _02713_;
  wire _02714_;
  wire _02715_;
  wire _02716_;
  wire _02717_;
  wire _02718_;
  wire _02719_;
  wire _02720_;
  wire _02721_;
  wire _02722_;
  wire _02723_;
  wire _02724_;
  wire _02725_;
  wire _02726_;
  wire _02727_;
  wire _02728_;
  wire _02729_;
  wire _02730_;
  wire _02731_;
  wire _02732_;
  wire _02733_;
  wire _02734_;
  wire _02735_;
  wire _02736_;
  wire _02737_;
  wire _02738_;
  wire _02739_;
  wire _02740_;
  wire _02741_;
  wire _02742_;
  wire _02743_;
  wire _02744_;
  wire _02745_;
  wire _02746_;
  wire _02747_;
  wire _02748_;
  wire _02749_;
  wire _02750_;
  wire _02751_;
  wire _02752_;
  wire _02753_;
  wire _02754_;
  wire _02755_;
  wire _02756_;
  wire _02757_;
  wire _02758_;
  wire _02759_;
  wire _02760_;
  wire _02761_;
  wire _02762_;
  wire _02763_;
  wire _02764_;
  wire _02765_;
  wire _02766_;
  wire _02767_;
  wire _02768_;
  wire _02769_;
  wire _02770_;
  wire _02771_;
  wire _02772_;
  wire _02773_;
  wire _02774_;
  wire _02775_;
  wire _02776_;
  wire _02777_;
  wire _02778_;
  wire _02779_;
  wire _02780_;
  wire _02781_;
  wire _02782_;
  wire _02783_;
  wire _02784_;
  wire _02785_;
  wire _02786_;
  wire _02787_;
  wire _02788_;
  wire _02789_;
  wire _02790_;
  wire _02791_;
  wire _02792_;
  wire _02793_;
  wire _02794_;
  wire _02795_;
  wire _02796_;
  wire _02797_;
  wire _02798_;
  wire _02799_;
  wire _02800_;
  wire _02801_;
  wire _02802_;
  wire _02803_;
  wire _02804_;
  wire _02805_;
  wire _02806_;
  wire _02807_;
  wire _02808_;
  wire _02809_;
  wire _02810_;
  wire _02811_;
  wire _02812_;
  wire _02813_;
  wire _02814_;
  wire _02815_;
  wire _02816_;
  wire _02817_;
  wire _02818_;
  wire _02819_;
  wire _02820_;
  wire _02821_;
  wire _02822_;
  wire _02823_;
  wire _02824_;
  wire _02825_;
  wire _02826_;
  wire _02827_;
  wire _02828_;
  wire _02829_;
  wire _02830_;
  wire _02831_;
  wire _02832_;
  wire _02833_;
  wire _02834_;
  wire _02835_;
  wire _02836_;
  wire _02837_;
  wire _02838_;
  wire _02839_;
  wire _02840_;
  wire _02841_;
  wire _02842_;
  wire _02843_;
  wire _02844_;
  wire _02845_;
  wire _02846_;
  wire _02847_;
  wire _02848_;
  wire _02849_;
  wire _02850_;
  wire _02851_;
  wire _02852_;
  wire _02853_;
  wire _02854_;
  wire _02855_;
  wire _02856_;
  wire _02857_;
  wire _02858_;
  wire _02859_;
  wire _02860_;
  wire _02861_;
  wire _02862_;
  wire _02863_;
  wire _02864_;
  wire _02865_;
  wire _02866_;
  wire _02867_;
  wire _02868_;
  wire _02869_;
  wire _02870_;
  wire _02871_;
  wire _02872_;
  wire _02873_;
  wire _02874_;
  wire _02875_;
  wire _02876_;
  wire _02877_;
  wire _02878_;
  wire _02879_;
  wire _02880_;
  wire _02881_;
  wire _02882_;
  wire _02883_;
  wire _02884_;
  wire _02885_;
  wire _02886_;
  wire _02887_;
  wire _02888_;
  wire _02889_;
  wire _02890_;
  wire _02891_;
  wire _02892_;
  wire _02893_;
  wire _02894_;
  wire _02895_;
  wire _02896_;
  wire _02897_;
  wire _02898_;
  wire _02899_;
  wire _02900_;
  wire _02901_;
  wire _02902_;
  wire _02903_;
  wire _02904_;
  wire _02905_;
  wire _02906_;
  wire _02907_;
  wire _02908_;
  wire _02909_;
  wire _02910_;
  wire _02911_;
  wire _02912_;
  wire _02913_;
  wire _02914_;
  wire _02915_;
  wire _02916_;
  wire _02917_;
  wire _02918_;
  wire _02919_;
  wire _02920_;
  wire _02921_;
  wire _02922_;
  wire _02923_;
  wire _02924_;
  wire _02925_;
  wire _02926_;
  wire _02927_;
  wire _02928_;
  wire _02929_;
  wire _02930_;
  wire _02931_;
  wire _02932_;
  wire _02933_;
  wire _02934_;
  wire _02935_;
  wire _02936_;
  wire _02937_;
  wire _02938_;
  wire _02939_;
  wire _02940_;
  wire _02941_;
  wire _02942_;
  wire _02943_;
  wire _02944_;
  wire _02945_;
  wire _02946_;
  wire _02947_;
  wire _02948_;
  wire _02949_;
  wire _02950_;
  wire _02951_;
  wire _02952_;
  wire _02953_;
  wire _02954_;
  wire _02955_;
  wire _02956_;
  wire _02957_;
  wire _02958_;
  wire _02959_;
  wire _02960_;
  wire _02961_;
  wire _02962_;
  wire _02963_;
  wire _02964_;
  wire _02965_;
  wire _02966_;
  wire _02967_;
  wire _02968_;
  wire _02969_;
  wire _02970_;
  wire _02971_;
  wire _02972_;
  wire _02973_;
  wire _02974_;
  wire _02975_;
  wire _02976_;
  wire _02977_;
  wire _02978_;
  wire _02979_;
  wire _02980_;
  wire _02981_;
  wire _02982_;
  wire _02983_;
  wire _02984_;
  wire _02985_;
  wire _02986_;
  wire _02987_;
  wire _02988_;
  wire _02989_;
  wire _02990_;
  wire _02991_;
  wire _02992_;
  wire _02993_;
  wire _02994_;
  wire _02995_;
  wire _02996_;
  wire _02997_;
  wire _02998_;
  wire _02999_;
  wire _03000_;
  wire _03001_;
  wire _03002_;
  wire _03003_;
  wire _03004_;
  wire _03005_;
  wire _03006_;
  wire _03007_;
  wire _03008_;
  wire _03009_;
  wire _03010_;
  wire _03011_;
  wire _03012_;
  wire _03013_;
  wire _03014_;
  wire _03015_;
  wire _03016_;
  wire _03017_;
  wire _03018_;
  wire _03019_;
  wire _03020_;
  wire _03021_;
  wire _03022_;
  wire _03023_;
  wire _03024_;
  wire _03025_;
  wire _03026_;
  wire _03027_;
  wire _03028_;
  wire _03029_;
  wire _03030_;
  wire _03031_;
  wire _03032_;
  wire _03033_;
  wire _03034_;
  wire _03035_;
  wire _03036_;
  wire _03037_;
  wire _03038_;
  wire _03039_;
  wire _03040_;
  wire _03041_;
  wire _03042_;
  wire _03043_;
  wire _03044_;
  wire _03045_;
  wire _03046_;
  wire _03047_;
  wire _03048_;
  wire _03049_;
  wire _03050_;
  wire _03051_;
  wire _03052_;
  wire _03053_;
  wire _03054_;
  wire _03055_;
  wire _03056_;
  wire _03057_;
  wire _03058_;
  wire _03059_;
  wire _03060_;
  wire _03061_;
  wire _03062_;
  wire _03063_;
  wire _03064_;
  wire _03065_;
  wire _03066_;
  wire _03067_;
  wire _03068_;
  wire _03069_;
  wire _03070_;
  wire _03071_;
  wire _03072_;
  wire _03073_;
  wire _03074_;
  wire _03075_;
  wire _03076_;
  wire _03077_;
  wire _03078_;
  wire _03079_;
  wire _03080_;
  wire _03081_;
  wire _03082_;
  wire _03083_;
  wire _03084_;
  wire _03085_;
  wire _03086_;
  wire _03087_;
  wire _03088_;
  wire _03089_;
  wire _03090_;
  wire _03091_;
  wire _03092_;
  wire _03093_;
  wire _03094_;
  wire _03095_;
  wire _03096_;
  wire _03097_;
  wire _03098_;
  wire _03099_;
  wire _03100_;
  wire _03101_;
  wire _03102_;
  wire _03103_;
  wire _03104_;
  wire _03105_;
  wire _03106_;
  wire _03107_;
  wire _03108_;
  wire _03109_;
  wire _03110_;
  wire _03111_;
  wire _03112_;
  wire _03113_;
  wire _03114_;
  wire _03115_;
  wire _03116_;
  wire _03117_;
  wire _03118_;
  wire _03119_;
  wire _03120_;
  wire _03121_;
  wire _03122_;
  wire _03123_;
  wire _03124_;
  wire _03125_;
  wire _03126_;
  wire _03127_;
  wire _03128_;
  wire _03129_;
  wire _03130_;
  wire _03131_;
  wire _03132_;
  wire _03133_;
  wire _03134_;
  wire _03135_;
  wire _03136_;
  wire _03137_;
  wire _03138_;
  wire _03139_;
  wire _03140_;
  wire _03141_;
  wire _03142_;
  wire _03143_;
  wire _03144_;
  wire _03145_;
  wire _03146_;
  wire _03147_;
  wire _03148_;
  wire _03149_;
  wire _03150_;
  wire _03151_;
  wire _03152_;
  wire _03153_;
  wire _03154_;
  wire _03155_;
  wire _03156_;
  wire _03157_;
  wire _03158_;
  wire _03159_;
  wire _03160_;
  wire _03161_;
  wire _03162_;
  wire _03163_;
  wire _03164_;
  wire _03165_;
  wire _03166_;
  wire _03167_;
  wire _03168_;
  wire _03169_;
  wire _03170_;
  wire _03171_;
  wire _03172_;
  wire _03173_;
  wire _03174_;
  wire _03175_;
  wire _03176_;
  wire _03177_;
  wire _03178_;
  wire _03179_;
  wire _03180_;
  wire _03181_;
  wire _03182_;
  wire _03183_;
  wire _03184_;
  wire _03185_;
  wire _03186_;
  wire _03187_;
  wire _03188_;
  wire _03189_;
  wire _03190_;
  wire _03191_;
  wire _03192_;
  wire _03193_;
  wire _03194_;
  wire _03195_;
  wire _03196_;
  wire _03197_;
  wire _03198_;
  wire _03199_;
  wire _03200_;
  wire _03201_;
  wire _03202_;
  wire _03203_;
  wire _03204_;
  wire _03205_;
  wire _03206_;
  wire _03207_;
  wire _03208_;
  wire _03209_;
  wire _03210_;
  wire _03211_;
  wire _03212_;
  wire _03213_;
  wire _03214_;
  wire _03215_;
  wire _03216_;
  wire _03217_;
  wire _03218_;
  wire _03219_;
  wire _03220_;
  wire _03221_;
  wire _03222_;
  wire _03223_;
  wire _03224_;
  wire _03225_;
  wire _03226_;
  wire _03227_;
  wire _03228_;
  wire _03229_;
  wire _03230_;
  wire _03231_;
  wire _03232_;
  wire _03233_;
  wire _03234_;
  wire _03235_;
  wire _03236_;
  wire _03237_;
  wire _03238_;
  wire _03239_;
  wire _03240_;
  wire _03241_;
  wire _03242_;
  wire _03243_;
  wire _03244_;
  wire _03245_;
  wire _03246_;
  wire _03247_;
  wire _03248_;
  wire _03249_;
  wire _03250_;
  wire _03251_;
  wire _03252_;
  wire _03253_;
  wire _03254_;
  wire _03255_;
  wire _03256_;
  wire _03257_;
  wire _03258_;
  wire _03259_;
  wire _03260_;
  wire _03261_;
  wire _03262_;
  wire _03263_;
  wire _03264_;
  wire _03265_;
  wire _03266_;
  wire _03267_;
  wire _03268_;
  wire _03269_;
  wire _03270_;
  wire _03271_;
  wire _03272_;
  wire _03273_;
  wire _03274_;
  wire _03275_;
  wire _03276_;
  wire _03277_;
  wire _03278_;
  wire _03279_;
  wire _03280_;
  wire _03281_;
  wire _03282_;
  wire _03283_;
  wire _03284_;
  wire _03285_;
  wire _03286_;
  wire _03287_;
  wire _03288_;
  wire _03289_;
  wire _03290_;
  wire _03291_;
  wire _03292_;
  wire _03293_;
  wire _03294_;
  wire _03295_;
  wire _03296_;
  wire _03297_;
  wire _03298_;
  wire _03299_;
  wire _03300_;
  wire _03301_;
  wire _03302_;
  wire _03303_;
  wire _03304_;
  wire _03305_;
  wire _03306_;
  wire _03307_;
  wire _03308_;
  wire _03309_;
  wire _03310_;
  wire _03311_;
  wire _03312_;
  wire _03313_;
  wire _03314_;
  wire _03315_;
  wire _03316_;
  wire _03317_;
  wire _03318_;
  wire _03319_;
  wire _03320_;
  wire _03321_;
  wire _03322_;
  wire _03323_;
  wire _03324_;
  wire _03325_;
  wire _03326_;
  wire _03327_;
  wire _03328_;
  wire _03329_;
  wire _03330_;
  wire _03331_;
  wire _03332_;
  wire _03333_;
  wire _03334_;
  wire _03335_;
  wire _03336_;
  wire _03337_;
  wire _03338_;
  wire _03339_;
  wire _03340_;
  wire _03341_;
  wire _03342_;
  wire _03343_;
  wire _03344_;
  wire _03345_;
  wire _03346_;
  wire _03347_;
  wire _03348_;
  wire _03349_;
  wire _03350_;
  wire _03351_;
  wire _03352_;
  wire _03353_;
  wire _03354_;
  wire _03355_;
  wire _03356_;
  wire _03357_;
  wire _03358_;
  wire _03359_;
  wire _03360_;
  wire _03361_;
  wire _03362_;
  wire _03363_;
  wire _03364_;
  wire _03365_;
  wire _03366_;
  wire _03367_;
  wire _03368_;
  wire _03369_;
  wire _03370_;
  wire _03371_;
  wire _03372_;
  wire _03373_;
  wire _03374_;
  wire _03375_;
  wire _03376_;
  wire _03377_;
  wire _03378_;
  wire _03379_;
  wire _03380_;
  wire _03381_;
  wire _03382_;
  wire _03383_;
  wire _03384_;
  wire _03385_;
  wire _03386_;
  wire _03387_;
  wire _03388_;
  wire _03389_;
  wire _03390_;
  wire _03391_;
  wire _03392_;
  wire _03393_;
  wire _03394_;
  wire _03395_;
  wire _03396_;
  wire _03397_;
  wire _03398_;
  wire _03399_;
  wire _03400_;
  wire _03401_;
  wire _03402_;
  wire _03403_;
  wire _03404_;
  wire _03405_;
  wire _03406_;
  wire _03407_;
  wire _03408_;
  wire _03409_;
  wire _03410_;
  wire _03411_;
  wire _03412_;
  wire _03413_;
  wire _03414_;
  wire _03415_;
  wire _03416_;
  wire _03417_;
  wire _03418_;
  wire _03419_;
  wire _03420_;
  wire _03421_;
  wire _03422_;
  wire _03423_;
  wire _03424_;
  wire _03425_;
  wire _03426_;
  wire _03427_;
  wire _03428_;
  wire _03429_;
  wire _03430_;
  wire _03431_;
  wire _03432_;
  wire _03433_;
  wire _03434_;
  wire _03435_;
  wire _03436_;
  wire _03437_;
  wire _03438_;
  wire _03439_;
  wire _03440_;
  wire _03441_;
  wire _03442_;
  wire _03443_;
  wire _03444_;
  wire _03445_;
  wire _03446_;
  wire _03447_;
  wire _03448_;
  wire _03449_;
  wire _03450_;
  wire _03451_;
  wire _03452_;
  wire _03453_;
  wire _03454_;
  wire _03455_;
  wire _03456_;
  wire _03457_;
  wire _03458_;
  wire _03459_;
  wire _03460_;
  wire _03461_;
  wire _03462_;
  wire _03463_;
  wire _03464_;
  wire _03465_;
  wire _03466_;
  wire _03467_;
  wire _03468_;
  wire _03469_;
  wire _03470_;
  wire _03471_;
  wire _03472_;
  wire _03473_;
  wire _03474_;
  wire _03475_;
  wire _03476_;
  wire _03477_;
  wire _03478_;
  wire _03479_;
  wire _03480_;
  wire _03481_;
  wire _03482_;
  wire _03483_;
  wire _03484_;
  wire _03485_;
  wire _03486_;
  wire _03487_;
  wire _03488_;
  wire _03489_;
  wire _03490_;
  wire _03491_;
  wire _03492_;
  wire _03493_;
  wire _03494_;
  wire _03495_;
  wire _03496_;
  wire _03497_;
  wire _03498_;
  wire _03499_;
  wire _03500_;
  wire _03501_;
  wire _03502_;
  wire _03503_;
  wire _03504_;
  wire _03505_;
  wire _03506_;
  wire _03507_;
  wire _03508_;
  wire _03509_;
  wire _03510_;
  wire _03511_;
  wire _03512_;
  wire _03513_;
  wire _03514_;
  wire _03515_;
  wire _03516_;
  wire _03517_;
  wire _03518_;
  wire _03519_;
  wire _03520_;
  wire _03521_;
  wire _03522_;
  wire _03523_;
  wire _03524_;
  wire _03525_;
  wire _03526_;
  wire _03527_;
  wire _03528_;
  wire _03529_;
  wire _03530_;
  wire _03531_;
  wire _03532_;
  wire _03533_;
  wire _03534_;
  wire _03535_;
  wire _03536_;
  wire _03537_;
  wire _03538_;
  wire _03539_;
  wire _03540_;
  wire _03541_;
  wire _03542_;
  wire _03543_;
  wire _03544_;
  wire _03545_;
  wire _03546_;
  wire _03547_;
  wire _03548_;
  wire _03549_;
  wire _03550_;
  wire _03551_;
  wire _03552_;
  wire _03553_;
  wire _03554_;
  wire _03555_;
  wire _03556_;
  wire _03557_;
  wire _03558_;
  wire _03559_;
  wire _03560_;
  wire _03561_;
  wire _03562_;
  wire _03563_;
  wire _03564_;
  wire _03565_;
  wire _03566_;
  wire _03567_;
  wire _03568_;
  wire _03569_;
  wire _03570_;
  wire _03571_;
  wire _03572_;
  wire _03573_;
  wire _03574_;
  wire _03575_;
  wire _03576_;
  wire _03577_;
  wire _03578_;
  wire _03579_;
  wire _03580_;
  wire _03581_;
  wire _03582_;
  wire _03583_;
  wire _03584_;
  wire _03585_;
  wire _03586_;
  wire _03587_;
  wire _03588_;
  wire _03589_;
  wire _03590_;
  wire _03591_;
  wire _03592_;
  wire _03593_;
  wire _03594_;
  wire _03595_;
  wire _03596_;
  wire _03597_;
  wire _03598_;
  wire _03599_;
  wire _03600_;
  wire _03601_;
  wire _03602_;
  wire _03603_;
  wire _03604_;
  wire _03605_;
  wire _03606_;
  wire _03607_;
  wire _03608_;
  wire _03609_;
  wire _03610_;
  wire _03611_;
  wire _03612_;
  wire _03613_;
  wire _03614_;
  wire _03615_;
  wire _03616_;
  wire _03617_;
  wire _03618_;
  wire _03619_;
  wire _03620_;
  wire _03621_;
  wire _03622_;
  wire _03623_;
  wire _03624_;
  wire _03625_;
  wire _03626_;
  wire _03627_;
  wire _03628_;
  wire _03629_;
  wire _03630_;
  wire _03631_;
  wire _03632_;
  wire _03633_;
  wire _03634_;
  wire _03635_;
  wire _03636_;
  wire _03637_;
  wire _03638_;
  wire _03639_;
  wire _03640_;
  wire _03641_;
  wire _03642_;
  wire _03643_;
  wire _03644_;
  wire _03645_;
  wire _03646_;
  wire _03647_;
  wire _03648_;
  wire _03649_;
  wire _03650_;
  wire _03651_;
  wire _03652_;
  wire _03653_;
  wire _03654_;
  wire _03655_;
  wire _03656_;
  wire _03657_;
  wire _03658_;
  wire _03659_;
  wire _03660_;
  wire _03661_;
  wire _03662_;
  wire _03663_;
  wire _03664_;
  wire _03665_;
  wire _03666_;
  wire _03667_;
  wire _03668_;
  wire _03669_;
  wire _03670_;
  wire _03671_;
  wire _03672_;
  wire _03673_;
  wire _03674_;
  wire _03675_;
  wire _03676_;
  wire _03677_;
  wire _03678_;
  wire _03679_;
  wire _03680_;
  wire _03681_;
  wire _03682_;
  wire _03683_;
  wire _03684_;
  wire _03685_;
  wire _03686_;
  wire _03687_;
  wire _03688_;
  wire _03689_;
  wire _03690_;
  wire _03691_;
  wire _03692_;
  wire _03693_;
  wire _03694_;
  wire _03695_;
  wire _03696_;
  wire _03697_;
  wire _03698_;
  wire _03699_;
  wire _03700_;
  wire _03701_;
  wire _03702_;
  wire _03703_;
  wire _03704_;
  wire _03705_;
  wire _03706_;
  wire _03707_;
  wire _03708_;
  wire _03709_;
  wire _03710_;
  wire _03711_;
  wire _03712_;
  wire _03713_;
  wire _03714_;
  wire _03715_;
  wire _03716_;
  wire _03717_;
  wire _03718_;
  wire _03719_;
  wire _03720_;
  wire _03721_;
  wire _03722_;
  wire _03723_;
  wire _03724_;
  wire _03725_;
  wire _03726_;
  wire _03727_;
  wire _03728_;
  wire _03729_;
  wire _03730_;
  wire _03731_;
  wire _03732_;
  wire _03733_;
  wire _03734_;
  wire _03735_;
  wire _03736_;
  wire _03737_;
  wire _03738_;
  wire _03739_;
  wire _03740_;
  wire _03741_;
  wire _03742_;
  wire _03743_;
  wire _03744_;
  wire _03745_;
  wire _03746_;
  wire _03747_;
  wire _03748_;
  wire _03749_;
  wire _03750_;
  wire _03751_;
  wire _03752_;
  wire _03753_;
  wire _03754_;
  wire _03755_;
  wire _03756_;
  wire _03757_;
  wire _03758_;
  wire _03759_;
  wire _03760_;
  wire _03761_;
  wire _03762_;
  wire _03763_;
  wire _03764_;
  wire _03765_;
  wire _03766_;
  wire _03767_;
  wire _03768_;
  wire _03769_;
  wire _03770_;
  wire _03771_;
  wire _03772_;
  wire _03773_;
  wire _03774_;
  wire _03775_;
  wire _03776_;
  wire _03777_;
  wire _03778_;
  wire _03779_;
  wire _03780_;
  wire _03781_;
  wire _03782_;
  wire _03783_;
  wire _03784_;
  wire _03785_;
  wire _03786_;
  wire _03787_;
  wire _03788_;
  wire _03789_;
  wire _03790_;
  wire _03791_;
  wire _03792_;
  wire _03793_;
  wire _03794_;
  wire _03795_;
  wire _03796_;
  wire _03797_;
  wire _03798_;
  wire _03799_;
  wire _03800_;
  wire _03801_;
  wire _03802_;
  wire _03803_;
  wire _03804_;
  wire _03805_;
  wire _03806_;
  wire _03807_;
  wire _03808_;
  wire _03809_;
  wire _03810_;
  wire _03811_;
  wire _03812_;
  wire _03813_;
  wire _03814_;
  wire _03815_;
  wire _03816_;
  wire _03817_;
  wire _03818_;
  wire _03819_;
  wire _03820_;
  wire _03821_;
  wire _03822_;
  wire _03823_;
  wire _03824_;
  wire _03825_;
  wire _03826_;
  wire _03827_;
  wire _03828_;
  wire _03829_;
  wire _03830_;
  wire _03831_;
  wire _03832_;
  wire _03833_;
  wire _03834_;
  wire _03835_;
  wire _03836_;
  wire _03837_;
  wire _03838_;
  wire _03839_;
  wire _03840_;
  wire _03841_;
  wire _03842_;
  wire _03843_;
  wire _03844_;
  wire _03845_;
  wire _03846_;
  wire _03847_;
  wire _03848_;
  wire _03849_;
  wire _03850_;
  wire _03851_;
  wire _03852_;
  wire _03853_;
  wire _03854_;
  wire _03855_;
  wire _03856_;
  wire _03857_;
  wire _03858_;
  wire _03859_;
  wire _03860_;
  wire _03861_;
  wire _03862_;
  wire _03863_;
  wire _03864_;
  wire _03865_;
  wire _03866_;
  wire _03867_;
  wire _03868_;
  wire _03869_;
  wire _03870_;
  wire _03871_;
  wire _03872_;
  wire _03873_;
  wire _03874_;
  wire _03875_;
  wire _03876_;
  wire _03877_;
  wire _03878_;
  wire _03879_;
  wire _03880_;
  wire _03881_;
  wire _03882_;
  wire _03883_;
  wire _03884_;
  wire _03885_;
  wire _03886_;
  wire _03887_;
  wire _03888_;
  wire _03889_;
  wire _03890_;
  wire _03891_;
  wire _03892_;
  wire _03893_;
  wire _03894_;
  wire _03895_;
  wire _03896_;
  wire _03897_;
  wire _03898_;
  wire _03899_;
  wire _03900_;
  wire _03901_;
  wire _03902_;
  wire _03903_;
  wire _03904_;
  wire _03905_;
  wire _03906_;
  wire _03907_;
  wire _03908_;
  wire _03909_;
  wire _03910_;
  wire _03911_;
  wire _03912_;
  wire _03913_;
  wire _03914_;
  wire _03915_;
  wire _03916_;
  wire _03917_;
  wire _03918_;
  wire _03919_;
  wire _03920_;
  wire _03921_;
  wire _03922_;
  wire _03923_;
  wire _03924_;
  wire _03925_;
  wire _03926_;
  wire _03927_;
  wire _03928_;
  wire _03929_;
  wire _03930_;
  wire _03931_;
  wire _03932_;
  wire _03933_;
  wire _03934_;
  wire _03935_;
  wire _03936_;
  wire _03937_;
  wire _03938_;
  wire _03939_;
  wire _03940_;
  wire _03941_;
  wire _03942_;
  wire _03943_;
  wire _03944_;
  wire _03945_;
  wire _03946_;
  wire _03947_;
  wire _03948_;
  wire _03949_;
  wire _03950_;
  wire _03951_;
  wire _03952_;
  wire _03953_;
  wire _03954_;
  wire _03955_;
  wire _03956_;
  wire _03957_;
  wire _03958_;
  wire _03959_;
  wire _03960_;
  wire _03961_;
  wire _03962_;
  wire _03963_;
  wire _03964_;
  wire _03965_;
  wire _03966_;
  wire _03967_;
  wire _03968_;
  wire _03969_;
  wire _03970_;
  wire _03971_;
  wire _03972_;
  wire _03973_;
  wire _03974_;
  wire _03975_;
  wire _03976_;
  wire _03977_;
  wire _03978_;
  wire _03979_;
  wire _03980_;
  wire _03981_;
  wire _03982_;
  wire _03983_;
  wire _03984_;
  wire _03985_;
  wire _03986_;
  wire _03987_;
  wire _03988_;
  wire _03989_;
  wire _03990_;
  wire _03991_;
  wire _03992_;
  wire _03993_;
  wire _03994_;
  wire _03995_;
  wire _03996_;
  wire _03997_;
  wire _03998_;
  wire _03999_;
  wire _04000_;
  wire _04001_;
  wire _04002_;
  wire _04003_;
  wire _04004_;
  wire _04005_;
  wire _04006_;
  wire _04007_;
  wire _04008_;
  wire _04009_;
  wire _04010_;
  wire _04011_;
  wire _04012_;
  wire _04013_;
  wire _04014_;
  wire _04015_;
  wire _04016_;
  wire _04017_;
  wire _04018_;
  wire _04019_;
  wire _04020_;
  wire _04021_;
  wire _04022_;
  wire _04023_;
  wire _04024_;
  wire _04025_;
  wire _04026_;
  wire _04027_;
  wire _04028_;
  wire _04029_;
  wire _04030_;
  wire _04031_;
  wire _04032_;
  wire _04033_;
  wire _04034_;
  wire _04035_;
  wire _04036_;
  wire _04037_;
  wire _04038_;
  wire _04039_;
  wire _04040_;
  wire _04041_;
  wire _04042_;
  wire _04043_;
  wire _04044_;
  wire _04045_;
  wire _04046_;
  wire _04047_;
  wire _04048_;
  wire _04049_;
  wire _04050_;
  wire _04051_;
  wire _04052_;
  wire _04053_;
  wire _04054_;
  wire _04055_;
  wire _04056_;
  wire _04057_;
  wire _04058_;
  wire _04059_;
  wire _04060_;
  wire _04061_;
  wire _04062_;
  wire _04063_;
  wire _04064_;
  wire _04065_;
  wire _04066_;
  wire _04067_;
  wire _04068_;
  wire _04069_;
  wire _04070_;
  wire _04071_;
  wire _04072_;
  wire _04073_;
  wire _04074_;
  wire _04075_;
  wire _04076_;
  wire _04077_;
  wire _04078_;
  wire _04079_;
  wire _04080_;
  wire _04081_;
  wire _04082_;
  wire _04083_;
  wire _04084_;
  wire _04085_;
  wire _04086_;
  wire _04087_;
  wire _04088_;
  wire _04089_;
  wire _04090_;
  wire _04091_;
  wire _04092_;
  wire _04093_;
  wire _04094_;
  wire _04095_;
  wire _04096_;
  wire _04097_;
  wire _04098_;
  wire _04099_;
  wire _04100_;
  wire _04101_;
  wire _04102_;
  wire _04103_;
  wire _04104_;
  wire _04105_;
  wire _04106_;
  wire _04107_;
  wire _04108_;
  wire _04109_;
  wire _04110_;
  wire _04111_;
  wire _04112_;
  wire _04113_;
  wire _04114_;
  wire _04115_;
  wire _04116_;
  wire _04117_;
  wire _04118_;
  wire _04119_;
  wire _04120_;
  wire _04121_;
  wire _04122_;
  wire _04123_;
  wire _04124_;
  wire _04125_;
  wire _04126_;
  wire _04127_;
  wire _04128_;
  wire _04129_;
  wire _04130_;
  wire _04131_;
  wire _04132_;
  wire _04133_;
  wire _04134_;
  wire _04135_;
  wire _04136_;
  wire _04137_;
  wire _04138_;
  wire _04139_;
  wire _04140_;
  wire _04141_;
  wire _04142_;
  wire _04143_;
  wire _04144_;
  wire _04145_;
  wire _04146_;
  wire _04147_;
  wire _04148_;
  wire _04149_;
  wire _04150_;
  wire _04151_;
  wire _04152_;
  wire _04153_;
  wire _04154_;
  wire _04155_;
  wire _04156_;
  wire _04157_;
  wire _04158_;
  wire _04159_;
  wire _04160_;
  wire _04161_;
  wire _04162_;
  wire _04163_;
  wire _04164_;
  wire _04165_;
  wire _04166_;
  wire _04167_;
  wire _04168_;
  wire _04169_;
  wire _04170_;
  wire _04171_;
  wire _04172_;
  wire _04173_;
  wire _04174_;
  wire _04175_;
  wire _04176_;
  wire _04177_;
  wire _04178_;
  wire _04179_;
  wire _04180_;
  wire _04181_;
  wire _04182_;
  wire _04183_;
  wire _04184_;
  wire _04185_;
  wire _04186_;
  wire _04187_;
  wire _04188_;
  wire _04189_;
  wire _04190_;
  wire _04191_;
  wire _04192_;
  wire _04193_;
  wire _04194_;
  wire _04195_;
  wire _04196_;
  wire _04197_;
  wire _04198_;
  wire _04199_;
  wire _04200_;
  wire _04201_;
  wire _04202_;
  wire _04203_;
  wire _04204_;
  wire _04205_;
  wire _04206_;
  wire _04207_;
  wire _04208_;
  wire _04209_;
  wire _04210_;
  wire _04211_;
  wire _04212_;
  wire _04213_;
  wire _04214_;
  wire _04215_;
  wire _04216_;
  wire _04217_;
  wire _04218_;
  wire _04219_;
  wire _04220_;
  wire _04221_;
  wire _04222_;
  wire _04223_;
  wire _04224_;
  wire _04225_;
  wire _04226_;
  wire _04227_;
  wire _04228_;
  wire _04229_;
  wire _04230_;
  wire _04231_;
  wire _04232_;
  wire _04233_;
  wire _04234_;
  wire _04235_;
  wire _04236_;
  wire _04237_;
  wire _04238_;
  wire _04239_;
  wire _04240_;
  wire _04241_;
  wire _04242_;
  wire _04243_;
  wire _04244_;
  wire _04245_;
  wire _04246_;
  wire _04247_;
  wire _04248_;
  wire _04249_;
  wire _04250_;
  wire _04251_;
  wire _04252_;
  wire _04253_;
  wire _04254_;
  wire _04255_;
  wire _04256_;
  wire _04257_;
  wire _04258_;
  wire _04259_;
  wire _04260_;
  wire _04261_;
  wire _04262_;
  wire _04263_;
  wire _04264_;
  wire _04265_;
  wire _04266_;
  wire _04267_;
  wire _04268_;
  wire _04269_;
  wire _04270_;
  wire _04271_;
  wire _04272_;
  wire _04273_;
  wire _04274_;
  wire _04275_;
  wire _04276_;
  wire _04277_;
  wire _04278_;
  wire _04279_;
  wire _04280_;
  wire _04281_;
  wire _04282_;
  wire _04283_;
  wire _04284_;
  wire _04285_;
  wire _04286_;
  wire _04287_;
  wire _04288_;
  wire _04289_;
  wire _04290_;
  wire _04291_;
  wire _04292_;
  wire _04293_;
  wire _04294_;
  wire _04295_;
  wire _04296_;
  wire _04297_;
  wire _04298_;
  wire _04299_;
  wire _04300_;
  wire _04301_;
  wire _04302_;
  wire _04303_;
  wire _04304_;
  wire _04305_;
  wire _04306_;
  wire _04307_;
  wire _04308_;
  wire _04309_;
  wire _04310_;
  wire _04311_;
  wire _04312_;
  wire _04313_;
  wire _04314_;
  wire _04315_;
  wire _04316_;
  wire _04317_;
  wire _04318_;
  wire _04319_;
  wire _04320_;
  wire _04321_;
  wire _04322_;
  wire _04323_;
  wire _04324_;
  wire _04325_;
  wire _04326_;
  wire _04327_;
  wire _04328_;
  wire _04329_;
  wire _04330_;
  wire _04331_;
  wire _04332_;
  wire _04333_;
  wire _04334_;
  wire _04335_;
  wire _04336_;
  wire _04337_;
  wire _04338_;
  wire _04339_;
  wire _04340_;
  wire _04341_;
  wire _04342_;
  wire _04343_;
  wire _04344_;
  wire _04345_;
  wire _04346_;
  wire _04347_;
  wire _04348_;
  wire _04349_;
  wire _04350_;
  wire _04351_;
  wire _04352_;
  wire _04353_;
  wire _04354_;
  wire _04355_;
  wire _04356_;
  wire _04357_;
  wire _04358_;
  wire _04359_;
  wire _04360_;
  wire _04361_;
  wire _04362_;
  wire _04363_;
  wire _04364_;
  wire _04365_;
  wire _04366_;
  wire _04367_;
  wire _04368_;
  wire _04369_;
  wire _04370_;
  wire _04371_;
  wire _04372_;
  wire _04373_;
  wire _04374_;
  wire _04375_;
  wire _04376_;
  wire _04377_;
  wire _04378_;
  wire _04379_;
  wire _04380_;
  wire _04381_;
  wire _04382_;
  wire _04383_;
  wire _04384_;
  wire _04385_;
  wire _04386_;
  wire _04387_;
  wire _04388_;
  wire _04389_;
  wire _04390_;
  wire _04391_;
  wire _04392_;
  wire _04393_;
  wire _04394_;
  wire _04395_;
  wire _04396_;
  wire _04397_;
  wire _04398_;
  wire _04399_;
  wire _04400_;
  wire _04401_;
  wire _04402_;
  wire _04403_;
  wire _04404_;
  wire _04405_;
  wire _04406_;
  wire _04407_;
  wire _04408_;
  wire _04409_;
  wire _04410_;
  wire _04411_;
  wire _04412_;
  wire _04413_;
  wire _04414_;
  wire _04415_;
  wire _04416_;
  wire _04417_;
  wire _04418_;
  wire _04419_;
  wire _04420_;
  wire _04421_;
  wire _04422_;
  wire _04423_;
  wire _04424_;
  wire _04425_;
  wire _04426_;
  wire _04427_;
  wire _04428_;
  wire _04429_;
  wire _04430_;
  wire _04431_;
  wire _04432_;
  wire _04433_;
  wire _04434_;
  wire _04435_;
  wire _04436_;
  wire _04437_;
  wire _04438_;
  wire _04439_;
  wire _04440_;
  wire _04441_;
  wire _04442_;
  wire _04443_;
  wire _04444_;
  wire _04445_;
  wire _04446_;
  wire _04447_;
  wire _04448_;
  wire _04449_;
  wire _04450_;
  wire _04451_;
  wire _04452_;
  wire _04453_;
  wire _04454_;
  wire _04455_;
  wire _04456_;
  wire _04457_;
  wire _04458_;
  wire _04459_;
  wire _04460_;
  wire _04461_;
  wire _04462_;
  wire _04463_;
  wire _04464_;
  wire _04465_;
  wire _04466_;
  wire _04467_;
  wire _04468_;
  wire _04469_;
  wire _04470_;
  wire _04471_;
  wire _04472_;
  wire _04473_;
  wire _04474_;
  wire _04475_;
  wire _04476_;
  wire _04477_;
  wire _04478_;
  wire _04479_;
  wire _04480_;
  wire _04481_;
  wire _04482_;
  wire _04483_;
  wire _04484_;
  wire _04485_;
  wire _04486_;
  wire _04487_;
  wire _04488_;
  wire _04489_;
  wire _04490_;
  wire _04491_;
  wire _04492_;
  wire _04493_;
  wire _04494_;
  wire _04495_;
  wire _04496_;
  wire _04497_;
  wire _04498_;
  wire _04499_;
  wire _04500_;
  wire _04501_;
  wire _04502_;
  wire _04503_;
  wire _04504_;
  wire _04505_;
  wire _04506_;
  wire _04507_;
  wire _04508_;
  wire _04509_;
  wire _04510_;
  wire _04511_;
  wire _04512_;
  wire _04513_;
  wire _04514_;
  wire _04515_;
  wire _04516_;
  wire _04517_;
  wire _04518_;
  wire _04519_;
  wire _04520_;
  wire _04521_;
  wire _04522_;
  wire _04523_;
  wire _04524_;
  wire _04525_;
  wire _04526_;
  wire _04527_;
  wire _04528_;
  wire _04529_;
  wire _04530_;
  wire _04531_;
  wire _04532_;
  wire _04533_;
  wire _04534_;
  wire _04535_;
  wire _04536_;
  wire _04537_;
  wire _04538_;
  wire _04539_;
  wire _04540_;
  wire _04541_;
  wire _04542_;
  wire _04543_;
  wire _04544_;
  wire _04545_;
  wire _04546_;
  wire _04547_;
  wire _04548_;
  wire _04549_;
  wire _04550_;
  wire _04551_;
  wire _04552_;
  wire _04553_;
  wire _04554_;
  wire _04555_;
  wire _04556_;
  wire _04557_;
  wire _04558_;
  wire _04559_;
  wire _04560_;
  wire _04561_;
  wire _04562_;
  wire _04563_;
  wire _04564_;
  wire _04565_;
  wire _04566_;
  wire _04567_;
  wire _04568_;
  wire _04569_;
  wire _04570_;
  wire _04571_;
  wire _04572_;
  wire _04573_;
  wire _04574_;
  wire _04575_;
  wire _04576_;
  wire _04577_;
  wire _04578_;
  wire _04579_;
  wire _04580_;
  wire _04581_;
  wire _04582_;
  wire _04583_;
  wire _04584_;
  wire _04585_;
  wire _04586_;
  wire _04587_;
  wire _04588_;
  wire _04589_;
  wire _04590_;
  wire _04591_;
  wire _04592_;
  wire _04593_;
  wire _04594_;
  wire _04595_;
  wire _04596_;
  wire _04597_;
  wire _04598_;
  wire _04599_;
  wire _04600_;
  wire _04601_;
  wire _04602_;
  wire _04603_;
  wire _04604_;
  wire _04605_;
  wire _04606_;
  wire _04607_;
  wire _04608_;
  wire _04609_;
  wire _04610_;
  wire _04611_;
  wire _04612_;
  wire _04613_;
  wire _04614_;
  wire _04615_;
  wire _04616_;
  wire _04617_;
  wire _04618_;
  wire _04619_;
  wire _04620_;
  wire _04621_;
  wire _04622_;
  wire _04623_;
  wire _04624_;
  wire _04625_;
  wire _04626_;
  wire _04627_;
  wire _04628_;
  wire _04629_;
  wire _04630_;
  wire _04631_;
  wire _04632_;
  wire _04633_;
  wire _04634_;
  wire _04635_;
  wire _04636_;
  wire _04637_;
  wire _04638_;
  wire _04639_;
  wire _04640_;
  wire _04641_;
  wire _04642_;
  wire _04643_;
  wire _04644_;
  wire _04645_;
  wire _04646_;
  wire _04647_;
  wire _04648_;
  wire _04649_;
  wire _04650_;
  wire _04651_;
  wire _04652_;
  wire _04653_;
  wire _04654_;
  wire _04655_;
  wire _04656_;
  wire _04657_;
  wire _04658_;
  wire _04659_;
  wire _04660_;
  wire _04661_;
  wire _04662_;
  wire _04663_;
  wire _04664_;
  wire _04665_;
  wire _04666_;
  wire _04667_;
  wire _04668_;
  wire _04669_;
  wire _04670_;
  wire _04671_;
  wire _04672_;
  wire _04673_;
  wire _04674_;
  wire _04675_;
  wire _04676_;
  wire _04677_;
  wire _04678_;
  wire _04679_;
  wire _04680_;
  wire _04681_;
  wire _04682_;
  wire _04683_;
  wire _04684_;
  wire _04685_;
  wire _04686_;
  wire _04687_;
  wire _04688_;
  wire _04689_;
  wire _04690_;
  wire _04691_;
  wire _04692_;
  wire _04693_;
  wire _04694_;
  wire _04695_;
  wire _04696_;
  wire _04697_;
  wire _04698_;
  wire _04699_;
  wire _04700_;
  wire _04701_;
  wire _04702_;
  wire _04703_;
  wire _04704_;
  wire _04705_;
  wire _04706_;
  wire _04707_;
  wire _04708_;
  wire _04709_;
  wire _04710_;
  wire _04711_;
  wire _04712_;
  wire _04713_;
  wire _04714_;
  wire _04715_;
  wire _04716_;
  wire _04717_;
  wire _04718_;
  wire _04719_;
  wire _04720_;
  wire _04721_;
  wire _04722_;
  wire _04723_;
  wire _04724_;
  wire _04725_;
  wire _04726_;
  wire _04727_;
  wire _04728_;
  wire _04729_;
  wire _04730_;
  wire _04731_;
  wire _04732_;
  wire _04733_;
  wire _04734_;
  wire _04735_;
  wire _04736_;
  wire _04737_;
  wire _04738_;
  wire _04739_;
  wire _04740_;
  wire _04741_;
  wire _04742_;
  wire _04743_;
  wire _04744_;
  wire _04745_;
  wire _04746_;
  wire _04747_;
  wire _04748_;
  wire _04749_;
  wire _04750_;
  wire _04751_;
  wire _04752_;
  wire _04753_;
  wire _04754_;
  wire _04755_;
  wire _04756_;
  wire _04757_;
  wire _04758_;
  wire _04759_;
  wire _04760_;
  wire _04761_;
  wire _04762_;
  wire _04763_;
  wire _04764_;
  wire _04765_;
  wire _04766_;
  wire _04767_;
  wire _04768_;
  wire _04769_;
  wire _04770_;
  wire _04771_;
  wire _04772_;
  wire _04773_;
  wire _04774_;
  wire _04775_;
  wire _04776_;
  wire _04777_;
  wire _04778_;
  wire _04779_;
  wire _04780_;
  wire _04781_;
  wire _04782_;
  wire _04783_;
  wire _04784_;
  wire _04785_;
  wire _04786_;
  wire _04787_;
  wire _04788_;
  wire _04789_;
  wire _04790_;
  wire _04791_;
  wire _04792_;
  wire _04793_;
  wire _04794_;
  wire _04795_;
  wire _04796_;
  wire _04797_;
  wire _04798_;
  wire _04799_;
  wire _04800_;
  wire _04801_;
  wire _04802_;
  wire _04803_;
  wire _04804_;
  wire _04805_;
  wire _04806_;
  wire _04807_;
  wire _04808_;
  wire _04809_;
  wire _04810_;
  wire _04811_;
  wire _04812_;
  wire _04813_;
  wire _04814_;
  wire _04815_;
  wire _04816_;
  wire _04817_;
  wire _04818_;
  wire _04819_;
  wire _04820_;
  wire _04821_;
  wire _04822_;
  wire _04823_;
  wire _04824_;
  wire _04825_;
  wire _04826_;
  wire _04827_;
  wire _04828_;
  wire _04829_;
  wire _04830_;
  wire _04831_;
  wire _04832_;
  wire _04833_;
  wire _04834_;
  wire _04835_;
  wire _04836_;
  wire _04837_;
  wire _04838_;
  wire _04839_;
  wire _04840_;
  wire _04841_;
  wire _04842_;
  wire _04843_;
  wire _04844_;
  wire _04845_;
  wire _04846_;
  wire _04847_;
  wire _04848_;
  wire _04849_;
  wire _04850_;
  wire _04851_;
  wire _04852_;
  wire _04853_;
  wire _04854_;
  wire _04855_;
  wire _04856_;
  wire _04857_;
  wire _04858_;
  wire _04859_;
  wire _04860_;
  wire _04861_;
  wire _04862_;
  wire _04863_;
  wire _04864_;
  wire _04865_;
  wire _04866_;
  wire _04867_;
  wire _04868_;
  wire _04869_;
  wire _04870_;
  wire _04871_;
  wire _04872_;
  wire _04873_;
  wire _04874_;
  wire _04875_;
  wire _04876_;
  wire _04877_;
  wire _04878_;
  wire _04879_;
  wire _04880_;
  wire _04881_;
  wire _04882_;
  wire _04883_;
  wire _04884_;
  wire _04885_;
  wire _04886_;
  wire _04887_;
  wire _04888_;
  wire _04889_;
  wire _04890_;
  wire _04891_;
  wire _04892_;
  wire _04893_;
  wire _04894_;
  wire _04895_;
  wire _04896_;
  wire _04897_;
  wire _04898_;
  wire _04899_;
  wire _04900_;
  wire _04901_;
  wire _04902_;
  wire _04903_;
  wire _04904_;
  wire _04905_;
  wire _04906_;
  wire _04907_;
  wire _04908_;
  wire _04909_;
  wire _04910_;
  wire _04911_;
  wire _04912_;
  wire _04913_;
  wire _04914_;
  wire _04915_;
  wire _04916_;
  wire _04917_;
  wire _04918_;
  wire _04919_;
  wire _04920_;
  wire _04921_;
  wire _04922_;
  wire _04923_;
  wire _04924_;
  wire _04925_;
  wire _04926_;
  wire _04927_;
  wire _04928_;
  wire _04929_;
  wire _04930_;
  wire _04931_;
  wire _04932_;
  wire _04933_;
  wire _04934_;
  wire _04935_;
  wire _04936_;
  wire _04937_;
  wire _04938_;
  wire _04939_;
  wire _04940_;
  wire _04941_;
  wire _04942_;
  wire _04943_;
  wire _04944_;
  wire _04945_;
  wire _04946_;
  wire _04947_;
  wire _04948_;
  wire _04949_;
  wire _04950_;
  wire _04951_;
  wire _04952_;
  wire _04953_;
  wire _04954_;
  wire _04955_;
  wire _04956_;
  wire _04957_;
  wire _04958_;
  wire _04959_;
  wire _04960_;
  wire _04961_;
  wire _04962_;
  wire _04963_;
  wire _04964_;
  wire _04965_;
  wire _04966_;
  wire _04967_;
  wire _04968_;
  wire _04969_;
  wire _04970_;
  wire _04971_;
  wire _04972_;
  wire _04973_;
  wire _04974_;
  wire _04975_;
  wire _04976_;
  wire _04977_;
  wire _04978_;
  wire _04979_;
  wire _04980_;
  wire _04981_;
  wire _04982_;
  wire _04983_;
  wire _04984_;
  wire _04985_;
  wire _04986_;
  wire _04987_;
  wire _04988_;
  wire _04989_;
  wire _04990_;
  wire _04991_;
  wire _04992_;
  wire _04993_;
  wire _04994_;
  wire _04995_;
  wire _04996_;
  wire _04997_;
  wire _04998_;
  wire _04999_;
  wire _05000_;
  wire _05001_;
  wire _05002_;
  wire _05003_;
  wire _05004_;
  wire _05005_;
  wire _05006_;
  wire _05007_;
  wire _05008_;
  wire _05009_;
  wire _05010_;
  wire _05011_;
  wire _05012_;
  wire _05013_;
  wire _05014_;
  wire _05015_;
  wire _05016_;
  wire _05017_;
  wire _05018_;
  wire _05019_;
  wire _05020_;
  wire _05021_;
  wire _05022_;
  wire _05023_;
  wire _05024_;
  wire _05025_;
  wire _05026_;
  wire _05027_;
  wire _05028_;
  wire _05029_;
  wire _05030_;
  wire _05031_;
  wire _05032_;
  wire _05033_;
  wire _05034_;
  wire _05035_;
  wire _05036_;
  wire _05037_;
  wire _05038_;
  wire _05039_;
  wire _05040_;
  wire _05041_;
  wire _05042_;
  wire _05043_;
  wire _05044_;
  wire _05045_;
  wire _05046_;
  wire _05047_;
  wire _05048_;
  wire _05049_;
  wire _05050_;
  wire _05051_;
  wire _05052_;
  wire _05053_;
  wire _05054_;
  wire _05055_;
  wire _05056_;
  wire _05057_;
  wire _05058_;
  wire _05059_;
  wire _05060_;
  wire _05061_;
  wire _05062_;
  wire _05063_;
  wire _05064_;
  wire _05065_;
  wire _05066_;
  wire _05067_;
  wire _05068_;
  wire _05069_;
  wire _05070_;
  wire _05071_;
  wire _05072_;
  wire _05073_;
  wire _05074_;
  wire _05075_;
  wire _05076_;
  wire _05077_;
  wire _05078_;
  wire _05079_;
  wire _05080_;
  wire _05081_;
  wire _05082_;
  wire _05083_;
  wire _05084_;
  wire _05085_;
  wire _05086_;
  wire _05087_;
  wire _05088_;
  wire _05089_;
  wire _05090_;
  wire _05091_;
  wire _05092_;
  wire _05093_;
  wire _05094_;
  wire _05095_;
  wire _05096_;
  wire _05097_;
  wire _05098_;
  wire _05099_;
  wire _05100_;
  wire _05101_;
  wire _05102_;
  wire _05103_;
  wire _05104_;
  wire _05105_;
  wire _05106_;
  wire _05107_;
  wire _05108_;
  wire _05109_;
  wire _05110_;
  wire _05111_;
  wire _05112_;
  wire _05113_;
  wire _05114_;
  wire _05115_;
  wire _05116_;
  wire _05117_;
  wire _05118_;
  wire _05119_;
  wire _05120_;
  wire _05121_;
  wire _05122_;
  wire _05123_;
  wire _05124_;
  wire _05125_;
  wire _05126_;
  wire _05127_;
  wire _05128_;
  wire _05129_;
  wire _05130_;
  wire _05131_;
  wire _05132_;
  wire _05133_;
  wire _05134_;
  wire _05135_;
  wire _05136_;
  wire _05137_;
  wire _05138_;
  wire _05139_;
  wire _05140_;
  wire _05141_;
  wire _05142_;
  wire _05143_;
  wire _05144_;
  wire _05145_;
  wire _05146_;
  wire _05147_;
  wire _05148_;
  wire _05149_;
  wire _05150_;
  wire _05151_;
  wire _05152_;
  wire _05153_;
  wire _05154_;
  wire _05155_;
  wire _05156_;
  wire _05157_;
  wire _05158_;
  wire _05159_;
  wire _05160_;
  wire _05161_;
  wire _05162_;
  wire _05163_;
  wire _05164_;
  wire _05165_;
  wire _05166_;
  wire _05167_;
  wire _05168_;
  wire _05169_;
  wire _05170_;
  wire _05171_;
  wire _05172_;
  wire _05173_;
  wire _05174_;
  wire _05175_;
  wire _05176_;
  wire _05177_;
  wire _05178_;
  wire _05179_;
  wire _05180_;
  wire _05181_;
  wire _05182_;
  wire _05183_;
  wire _05184_;
  wire _05185_;
  wire _05186_;
  wire _05187_;
  wire _05188_;
  wire _05189_;
  wire _05190_;
  wire _05191_;
  wire _05192_;
  wire _05193_;
  wire _05194_;
  wire _05195_;
  wire _05196_;
  wire _05197_;
  wire _05198_;
  wire _05199_;
  wire _05200_;
  wire _05201_;
  wire _05202_;
  wire _05203_;
  wire _05204_;
  wire _05205_;
  wire _05206_;
  wire _05207_;
  wire _05208_;
  wire _05209_;
  wire _05210_;
  wire _05211_;
  wire _05212_;
  wire _05213_;
  wire _05214_;
  wire _05215_;
  wire _05216_;
  wire _05217_;
  wire _05218_;
  wire _05219_;
  wire _05220_;
  wire _05221_;
  wire _05222_;
  wire _05223_;
  wire _05224_;
  wire _05225_;
  wire _05226_;
  wire _05227_;
  wire _05228_;
  wire _05229_;
  wire _05230_;
  wire _05231_;
  wire _05232_;
  wire _05233_;
  wire _05234_;
  wire _05235_;
  wire _05236_;
  wire _05237_;
  wire _05238_;
  wire _05239_;
  wire _05240_;
  wire _05241_;
  wire _05242_;
  wire _05243_;
  wire _05244_;
  wire _05245_;
  wire _05246_;
  wire _05247_;
  wire _05248_;
  wire _05249_;
  wire _05250_;
  wire _05251_;
  wire _05252_;
  wire _05253_;
  wire _05254_;
  wire _05255_;
  wire _05256_;
  wire _05257_;
  wire _05258_;
  wire _05259_;
  wire _05260_;
  wire _05261_;
  wire _05262_;
  wire _05263_;
  wire _05264_;
  wire _05265_;
  wire _05266_;
  wire _05267_;
  wire _05268_;
  wire _05269_;
  wire _05270_;
  wire _05271_;
  wire _05272_;
  wire _05273_;
  wire _05274_;
  wire _05275_;
  wire _05276_;
  wire _05277_;
  wire _05278_;
  wire _05279_;
  wire _05280_;
  wire _05281_;
  wire _05282_;
  wire _05283_;
  wire _05284_;
  wire _05285_;
  wire _05286_;
  wire _05287_;
  wire _05288_;
  wire _05289_;
  wire _05290_;
  wire _05291_;
  wire _05292_;
  wire _05293_;
  wire _05294_;
  wire _05295_;
  wire _05296_;
  wire _05297_;
  wire _05298_;
  wire _05299_;
  wire _05300_;
  wire _05301_;
  wire _05302_;
  wire _05303_;
  wire _05304_;
  wire _05305_;
  wire _05306_;
  wire _05307_;
  wire _05308_;
  wire _05309_;
  wire _05310_;
  wire _05311_;
  wire _05312_;
  wire _05313_;
  wire _05314_;
  wire _05315_;
  wire _05316_;
  wire _05317_;
  wire _05318_;
  wire _05319_;
  wire _05320_;
  wire _05321_;
  wire _05322_;
  wire _05323_;
  wire _05324_;
  wire _05325_;
  wire _05326_;
  wire _05327_;
  wire _05328_;
  wire _05329_;
  wire _05330_;
  wire _05331_;
  wire _05332_;
  wire _05333_;
  wire _05334_;
  wire _05335_;
  wire _05336_;
  wire _05337_;
  wire _05338_;
  wire _05339_;
  wire _05340_;
  wire _05341_;
  wire _05342_;
  wire _05343_;
  wire _05344_;
  wire _05345_;
  wire _05346_;
  wire _05347_;
  wire _05348_;
  wire _05349_;
  wire _05350_;
  wire _05351_;
  wire _05352_;
  wire _05353_;
  wire _05354_;
  wire _05355_;
  wire _05356_;
  wire _05357_;
  wire _05358_;
  wire _05359_;
  wire _05360_;
  wire _05361_;
  wire _05362_;
  wire _05363_;
  wire _05364_;
  wire _05365_;
  wire _05366_;
  wire _05367_;
  wire _05368_;
  wire _05369_;
  wire _05370_;
  wire _05371_;
  wire _05372_;
  wire _05373_;
  wire _05374_;
  wire _05375_;
  wire _05376_;
  wire _05377_;
  wire _05378_;
  wire _05379_;
  wire _05380_;
  wire _05381_;
  wire _05382_;
  wire _05383_;
  wire _05384_;
  wire _05385_;
  wire _05386_;
  wire _05387_;
  wire _05388_;
  wire _05389_;
  wire _05390_;
  wire _05391_;
  wire _05392_;
  wire _05393_;
  wire _05394_;
  wire _05395_;
  wire _05396_;
  wire _05397_;
  wire _05398_;
  wire _05399_;
  wire _05400_;
  wire _05401_;
  wire _05402_;
  wire _05403_;
  wire _05404_;
  wire _05405_;
  wire _05406_;
  wire _05407_;
  wire _05408_;
  wire _05409_;
  wire _05410_;
  wire _05411_;
  wire _05412_;
  wire _05413_;
  wire _05414_;
  wire _05415_;
  wire _05416_;
  wire _05417_;
  wire _05418_;
  wire _05419_;
  wire _05420_;
  wire _05421_;
  wire _05422_;
  wire _05423_;
  wire _05424_;
  wire _05425_;
  wire _05426_;
  wire _05427_;
  wire _05428_;
  wire _05429_;
  wire _05430_;
  wire _05431_;
  wire _05432_;
  wire _05433_;
  wire _05434_;
  wire _05435_;
  wire _05436_;
  wire _05437_;
  wire _05438_;
  wire _05439_;
  wire _05440_;
  wire _05441_;
  wire _05442_;
  wire _05443_;
  wire _05444_;
  wire _05445_;
  wire _05446_;
  wire _05447_;
  wire _05448_;
  wire _05449_;
  wire _05450_;
  wire _05451_;
  wire _05452_;
  wire _05453_;
  wire _05454_;
  wire _05455_;
  wire _05456_;
  wire _05457_;
  wire _05458_;
  wire _05459_;
  wire _05460_;
  wire _05461_;
  wire _05462_;
  wire _05463_;
  wire _05464_;
  wire _05465_;
  wire _05466_;
  wire _05467_;
  wire _05468_;
  wire _05469_;
  wire _05470_;
  wire _05471_;
  wire _05472_;
  wire _05473_;
  wire _05474_;
  wire _05475_;
  wire _05476_;
  wire _05477_;
  wire _05478_;
  wire _05479_;
  wire _05480_;
  wire _05481_;
  wire _05482_;
  wire _05483_;
  wire _05484_;
  wire _05485_;
  wire _05486_;
  wire _05487_;
  wire _05488_;
  wire _05489_;
  wire _05490_;
  wire _05491_;
  wire _05492_;
  wire _05493_;
  wire _05494_;
  wire _05495_;
  wire _05496_;
  wire _05497_;
  wire _05498_;
  wire _05499_;
  wire _05500_;
  wire _05501_;
  wire _05502_;
  wire _05503_;
  wire _05504_;
  wire _05505_;
  wire _05506_;
  wire _05507_;
  wire _05508_;
  wire _05509_;
  wire _05510_;
  wire _05511_;
  wire _05512_;
  wire _05513_;
  wire _05514_;
  wire _05515_;
  wire _05516_;
  wire _05517_;
  wire _05518_;
  wire _05519_;
  wire _05520_;
  wire _05521_;
  wire _05522_;
  wire _05523_;
  wire _05524_;
  wire _05525_;
  wire _05526_;
  wire _05527_;
  wire _05528_;
  wire _05529_;
  wire _05530_;
  wire _05531_;
  wire _05532_;
  wire _05533_;
  wire _05534_;
  wire _05535_;
  wire _05536_;
  wire _05537_;
  wire _05538_;
  wire _05539_;
  wire _05540_;
  wire _05541_;
  wire _05542_;
  wire _05543_;
  wire _05544_;
  wire _05545_;
  wire _05546_;
  wire _05547_;
  wire _05548_;
  wire _05549_;
  wire _05550_;
  wire _05551_;
  wire _05552_;
  wire _05553_;
  wire _05554_;
  wire _05555_;
  wire _05556_;
  wire _05557_;
  wire _05558_;
  wire _05559_;
  wire _05560_;
  wire _05561_;
  wire _05562_;
  wire _05563_;
  wire _05564_;
  wire _05565_;
  wire _05566_;
  wire _05567_;
  wire _05568_;
  wire _05569_;
  wire _05570_;
  wire _05571_;
  wire _05572_;
  wire _05573_;
  wire _05574_;
  wire _05575_;
  wire _05576_;
  wire _05577_;
  wire _05578_;
  wire _05579_;
  wire _05580_;
  wire _05581_;
  wire _05582_;
  wire _05583_;
  wire _05584_;
  wire _05585_;
  wire _05586_;
  wire _05587_;
  wire _05588_;
  wire _05589_;
  wire _05590_;
  wire _05591_;
  wire _05592_;
  wire _05593_;
  wire _05594_;
  wire _05595_;
  wire _05596_;
  wire _05597_;
  wire _05598_;
  wire _05599_;
  wire _05600_;
  wire _05601_;
  wire _05602_;
  wire _05603_;
  wire _05604_;
  wire _05605_;
  wire _05606_;
  wire _05607_;
  wire _05608_;
  wire _05609_;
  wire _05610_;
  wire _05611_;
  wire _05612_;
  wire _05613_;
  wire _05614_;
  wire _05615_;
  wire _05616_;
  wire _05617_;
  wire _05618_;
  wire _05619_;
  wire _05620_;
  wire _05621_;
  wire _05622_;
  wire _05623_;
  wire _05624_;
  wire _05625_;
  wire _05626_;
  wire _05627_;
  wire _05628_;
  wire _05629_;
  wire _05630_;
  wire _05631_;
  wire _05632_;
  wire _05633_;
  wire _05634_;
  wire _05635_;
  wire _05636_;
  wire _05637_;
  wire _05638_;
  wire _05639_;
  wire _05640_;
  wire _05641_;
  wire _05642_;
  wire _05643_;
  wire _05644_;
  wire _05645_;
  wire _05646_;
  wire _05647_;
  wire _05648_;
  wire _05649_;
  wire _05650_;
  wire _05651_;
  wire _05652_;
  wire _05653_;
  wire _05654_;
  wire _05655_;
  wire _05656_;
  wire _05657_;
  wire _05658_;
  wire _05659_;
  wire _05660_;
  wire _05661_;
  wire _05662_;
  wire _05663_;
  wire _05664_;
  wire _05665_;
  wire _05666_;
  wire _05667_;
  wire _05668_;
  wire _05669_;
  wire _05670_;
  wire _05671_;
  wire _05672_;
  wire _05673_;
  wire _05674_;
  wire _05675_;
  wire _05676_;
  wire _05677_;
  wire _05678_;
  wire _05679_;
  wire _05680_;
  wire _05681_;
  wire _05682_;
  wire _05683_;
  wire _05684_;
  wire _05685_;
  wire _05686_;
  wire _05687_;
  wire _05688_;
  wire _05689_;
  wire _05690_;
  wire _05691_;
  wire _05692_;
  wire _05693_;
  wire _05694_;
  wire _05695_;
  wire _05696_;
  wire _05697_;
  wire _05698_;
  wire _05699_;
  wire _05700_;
  wire _05701_;
  wire _05702_;
  wire _05703_;
  wire _05704_;
  wire _05705_;
  wire _05706_;
  wire _05707_;
  wire _05708_;
  wire _05709_;
  wire _05710_;
  wire _05711_;
  wire _05712_;
  wire _05713_;
  wire _05714_;
  wire _05715_;
  wire _05716_;
  wire _05717_;
  wire _05718_;
  wire _05719_;
  wire _05720_;
  wire _05721_;
  wire _05722_;
  wire _05723_;
  wire _05724_;
  wire _05725_;
  wire _05726_;
  wire _05727_;
  wire _05728_;
  wire _05729_;
  wire _05730_;
  wire _05731_;
  wire _05732_;
  wire _05733_;
  wire _05734_;
  wire _05735_;
  wire _05736_;
  wire _05737_;
  wire _05738_;
  wire _05739_;
  wire _05740_;
  wire _05741_;
  wire _05742_;
  wire _05743_;
  wire _05744_;
  wire _05745_;
  wire _05746_;
  wire _05747_;
  wire _05748_;
  wire _05749_;
  wire _05750_;
  wire _05751_;
  wire _05752_;
  wire _05753_;
  wire _05754_;
  wire _05755_;
  wire _05756_;
  wire _05757_;
  wire _05758_;
  wire _05759_;
  wire _05760_;
  wire _05761_;
  wire _05762_;
  wire _05763_;
  wire _05764_;
  wire _05765_;
  wire _05766_;
  wire _05767_;
  wire _05768_;
  wire _05769_;
  wire _05770_;
  wire _05771_;
  wire _05772_;
  wire _05773_;
  wire _05774_;
  wire _05775_;
  wire _05776_;
  wire _05777_;
  wire _05778_;
  wire _05779_;
  wire _05780_;
  wire _05781_;
  wire _05782_;
  wire _05783_;
  wire _05784_;
  wire _05785_;
  wire _05786_;
  wire _05787_;
  wire _05788_;
  wire _05789_;
  wire _05790_;
  wire _05791_;
  wire _05792_;
  wire _05793_;
  wire _05794_;
  wire _05795_;
  wire _05796_;
  wire _05797_;
  wire _05798_;
  wire _05799_;
  wire _05800_;
  wire _05801_;
  wire _05802_;
  wire _05803_;
  wire _05804_;
  wire _05805_;
  wire _05806_;
  wire _05807_;
  wire _05808_;
  wire _05809_;
  wire _05810_;
  wire _05811_;
  wire _05812_;
  wire _05813_;
  wire _05814_;
  wire _05815_;
  wire _05816_;
  wire _05817_;
  wire _05818_;
  wire _05819_;
  wire _05820_;
  wire _05821_;
  wire _05822_;
  wire _05823_;
  wire _05824_;
  wire _05825_;
  wire _05826_;
  wire _05827_;
  wire _05828_;
  wire _05829_;
  wire _05830_;
  wire _05831_;
  wire _05832_;
  wire _05833_;
  wire _05834_;
  wire _05835_;
  wire _05836_;
  wire _05837_;
  wire _05838_;
  wire _05839_;
  wire _05840_;
  wire _05841_;
  wire _05842_;
  wire _05843_;
  wire _05844_;
  wire _05845_;
  wire _05846_;
  wire _05847_;
  wire _05848_;
  wire _05849_;
  wire _05850_;
  wire _05851_;
  wire _05852_;
  wire _05853_;
  wire _05854_;
  wire _05855_;
  wire _05856_;
  wire _05857_;
  wire _05858_;
  wire _05859_;
  wire _05860_;
  wire _05861_;
  wire _05862_;
  wire _05863_;
  wire _05864_;
  wire _05865_;
  wire _05866_;
  wire _05867_;
  wire _05868_;
  wire _05869_;
  wire _05870_;
  wire _05871_;
  wire _05872_;
  wire _05873_;
  wire _05874_;
  wire _05875_;
  wire _05876_;
  wire _05877_;
  wire _05878_;
  wire _05879_;
  wire _05880_;
  wire _05881_;
  wire _05882_;
  wire _05883_;
  wire _05884_;
  wire _05885_;
  wire _05886_;
  wire _05887_;
  wire _05888_;
  wire _05889_;
  wire _05890_;
  wire _05891_;
  wire _05892_;
  wire _05893_;
  wire _05894_;
  wire _05895_;
  wire _05896_;
  wire _05897_;
  wire _05898_;
  wire _05899_;
  wire _05900_;
  wire _05901_;
  wire _05902_;
  wire _05903_;
  wire _05904_;
  wire _05905_;
  wire _05906_;
  wire _05907_;
  wire _05908_;
  wire _05909_;
  wire _05910_;
  wire _05911_;
  wire _05912_;
  wire _05913_;
  wire _05914_;
  wire _05915_;
  wire _05916_;
  wire _05917_;
  wire _05918_;
  wire _05919_;
  wire _05920_;
  wire _05921_;
  wire _05922_;
  wire _05923_;
  wire _05924_;
  wire _05925_;
  wire _05926_;
  wire _05927_;
  wire _05928_;
  wire _05929_;
  wire _05930_;
  wire _05931_;
  wire _05932_;
  wire _05933_;
  wire _05934_;
  wire _05935_;
  wire _05936_;
  wire _05937_;
  wire _05938_;
  wire _05939_;
  wire _05940_;
  wire _05941_;
  wire _05942_;
  wire _05943_;
  wire _05944_;
  wire _05945_;
  wire _05946_;
  wire _05947_;
  wire _05948_;
  wire _05949_;
  wire _05950_;
  wire _05951_;
  wire _05952_;
  wire _05953_;
  wire _05954_;
  wire _05955_;
  wire _05956_;
  wire _05957_;
  wire _05958_;
  wire _05959_;
  wire _05960_;
  wire _05961_;
  wire _05962_;
  wire _05963_;
  wire _05964_;
  wire _05965_;
  wire _05966_;
  wire _05967_;
  wire _05968_;
  wire _05969_;
  wire _05970_;
  wire _05971_;
  wire _05972_;
  wire _05973_;
  wire _05974_;
  wire _05975_;
  wire _05976_;
  wire _05977_;
  wire _05978_;
  wire _05979_;
  wire _05980_;
  wire _05981_;
  wire _05982_;
  wire _05983_;
  wire _05984_;
  wire _05985_;
  wire _05986_;
  wire _05987_;
  wire _05988_;
  wire _05989_;
  wire _05990_;
  wire _05991_;
  wire _05992_;
  wire _05993_;
  wire _05994_;
  wire _05995_;
  wire _05996_;
  wire _05997_;
  wire _05998_;
  wire _05999_;
  wire _06000_;
  wire _06001_;
  wire _06002_;
  wire _06003_;
  wire _06004_;
  wire _06005_;
  wire _06006_;
  wire _06007_;
  wire _06008_;
  wire _06009_;
  wire _06010_;
  wire _06011_;
  wire _06012_;
  wire _06013_;
  wire _06014_;
  wire _06015_;
  wire _06016_;
  wire _06017_;
  wire _06018_;
  wire _06019_;
  wire _06020_;
  wire _06021_;
  wire _06022_;
  wire _06023_;
  wire _06024_;
  wire _06025_;
  wire _06026_;
  wire _06027_;
  wire _06028_;
  wire _06029_;
  wire _06030_;
  wire _06031_;
  wire _06032_;
  wire _06033_;
  wire _06034_;
  wire _06035_;
  wire _06036_;
  wire _06037_;
  wire _06038_;
  wire _06039_;
  wire _06040_;
  wire _06041_;
  wire _06042_;
  wire _06043_;
  wire _06044_;
  wire _06045_;
  wire _06046_;
  wire _06047_;
  wire _06048_;
  wire _06049_;
  wire _06050_;
  wire _06051_;
  wire _06052_;
  wire _06053_;
  wire _06054_;
  wire _06055_;
  wire _06056_;
  wire _06057_;
  wire _06058_;
  wire _06059_;
  wire _06060_;
  wire _06061_;
  wire _06062_;
  wire _06063_;
  wire _06064_;
  wire _06065_;
  wire _06066_;
  wire _06067_;
  wire _06068_;
  wire _06069_;
  wire _06070_;
  wire _06071_;
  wire _06072_;
  wire _06073_;
  wire _06074_;
  wire _06075_;
  wire _06076_;
  wire _06077_;
  wire _06078_;
  wire _06079_;
  wire _06080_;
  wire _06081_;
  wire _06082_;
  wire _06083_;
  wire _06084_;
  wire _06085_;
  wire _06086_;
  wire _06087_;
  wire _06088_;
  wire _06089_;
  wire _06090_;
  wire _06091_;
  wire _06092_;
  wire _06093_;
  wire _06094_;
  wire _06095_;
  wire _06096_;
  wire _06097_;
  wire _06098_;
  wire _06099_;
  wire _06100_;
  wire _06101_;
  wire _06102_;
  wire _06103_;
  wire _06104_;
  wire _06105_;
  wire _06106_;
  wire _06107_;
  wire _06108_;
  wire _06109_;
  wire _06110_;
  wire _06111_;
  wire _06112_;
  wire _06113_;
  wire _06114_;
  wire _06115_;
  wire _06116_;
  wire _06117_;
  wire _06118_;
  wire _06119_;
  wire _06120_;
  wire _06121_;
  wire _06122_;
  wire _06123_;
  wire _06124_;
  wire _06125_;
  wire _06126_;
  wire _06127_;
  wire _06128_;
  wire _06129_;
  wire _06130_;
  wire _06131_;
  wire _06132_;
  wire _06133_;
  wire _06134_;
  wire _06135_;
  wire _06136_;
  wire _06137_;
  wire _06138_;
  wire _06139_;
  wire _06140_;
  wire _06141_;
  wire _06142_;
  wire _06143_;
  wire _06144_;
  wire _06145_;
  wire _06146_;
  wire _06147_;
  wire _06148_;
  wire _06149_;
  wire _06150_;
  wire _06151_;
  wire _06152_;
  wire _06153_;
  wire _06154_;
  wire _06155_;
  wire _06156_;
  wire _06157_;
  wire _06158_;
  wire _06159_;
  wire _06160_;
  wire _06161_;
  wire _06162_;
  wire _06163_;
  wire _06164_;
  wire _06165_;
  wire _06166_;
  wire _06167_;
  wire _06168_;
  wire _06169_;
  wire _06170_;
  wire _06171_;
  wire _06172_;
  wire _06173_;
  wire _06174_;
  wire _06175_;
  wire _06176_;
  wire _06177_;
  wire _06178_;
  wire _06179_;
  wire _06180_;
  wire _06181_;
  wire _06182_;
  wire _06183_;
  wire _06184_;
  wire _06185_;
  wire _06186_;
  wire _06187_;
  wire _06188_;
  wire _06189_;
  wire _06190_;
  wire _06191_;
  wire _06192_;
  wire _06193_;
  wire _06194_;
  wire _06195_;
  wire _06196_;
  wire _06197_;
  wire _06198_;
  wire _06199_;
  wire _06200_;
  wire _06201_;
  wire _06202_;
  wire _06203_;
  wire _06204_;
  wire _06205_;
  wire _06206_;
  wire _06207_;
  wire _06208_;
  wire _06209_;
  wire _06210_;
  wire _06211_;
  wire _06212_;
  wire _06213_;
  wire _06214_;
  wire _06215_;
  wire _06216_;
  wire _06217_;
  wire _06218_;
  wire _06219_;
  wire _06220_;
  wire _06221_;
  wire _06222_;
  wire _06223_;
  wire _06224_;
  wire _06225_;
  wire _06226_;
  wire _06227_;
  wire _06228_;
  wire _06229_;
  wire _06230_;
  wire _06231_;
  wire _06232_;
  wire _06233_;
  wire _06234_;
  wire _06235_;
  wire _06236_;
  wire _06237_;
  wire _06238_;
  wire _06239_;
  wire _06240_;
  wire _06241_;
  wire _06242_;
  wire _06243_;
  wire _06244_;
  wire _06245_;
  wire _06246_;
  wire _06247_;
  wire _06248_;
  wire _06249_;
  wire _06250_;
  wire _06251_;
  wire _06252_;
  wire _06253_;
  wire _06254_;
  wire _06255_;
  wire _06256_;
  wire _06257_;
  wire _06258_;
  wire _06259_;
  wire _06260_;
  wire _06261_;
  wire _06262_;
  wire _06263_;
  wire _06264_;
  wire _06265_;
  wire _06266_;
  wire _06267_;
  wire _06268_;
  wire _06269_;
  wire _06270_;
  wire _06271_;
  wire _06272_;
  wire _06273_;
  wire _06274_;
  wire _06275_;
  wire _06276_;
  wire _06277_;
  wire _06278_;
  wire _06279_;
  wire _06280_;
  wire _06281_;
  wire _06282_;
  wire _06283_;
  wire _06284_;
  wire _06285_;
  wire _06286_;
  wire _06287_;
  wire _06288_;
  wire _06289_;
  wire _06290_;
  wire _06291_;
  wire _06292_;
  wire _06293_;
  wire _06294_;
  wire _06295_;
  wire _06296_;
  wire _06297_;
  wire _06298_;
  wire _06299_;
  wire _06300_;
  wire _06301_;
  wire _06302_;
  wire _06303_;
  wire _06304_;
  wire _06305_;
  wire _06306_;
  wire _06307_;
  wire _06308_;
  wire _06309_;
  wire _06310_;
  wire _06311_;
  wire _06312_;
  wire _06313_;
  wire _06314_;
  wire _06315_;
  wire _06316_;
  wire _06317_;
  wire _06318_;
  wire _06319_;
  wire _06320_;
  wire _06321_;
  wire _06322_;
  wire _06323_;
  wire _06324_;
  wire _06325_;
  wire _06326_;
  wire _06327_;
  wire _06328_;
  wire _06329_;
  wire _06330_;
  wire _06331_;
  wire _06332_;
  wire _06333_;
  wire _06334_;
  wire _06335_;
  wire _06336_;
  wire _06337_;
  wire _06338_;
  wire _06339_;
  wire _06340_;
  wire _06341_;
  wire _06342_;
  wire _06343_;
  wire _06344_;
  wire _06345_;
  wire _06346_;
  wire _06347_;
  wire _06348_;
  wire _06349_;
  wire _06350_;
  wire _06351_;
  wire _06352_;
  wire _06353_;
  wire _06354_;
  wire _06355_;
  wire _06356_;
  wire _06357_;
  wire _06358_;
  wire _06359_;
  wire _06360_;
  wire _06361_;
  wire _06362_;
  wire _06363_;
  wire _06364_;
  wire _06365_;
  wire _06366_;
  wire _06367_;
  wire _06368_;
  wire _06369_;
  wire _06370_;
  wire _06371_;
  wire _06372_;
  wire _06373_;
  wire _06374_;
  wire _06375_;
  wire _06376_;
  wire _06377_;
  wire _06378_;
  wire _06379_;
  wire _06380_;
  wire _06381_;
  wire _06382_;
  wire _06383_;
  wire _06384_;
  wire _06385_;
  wire _06386_;
  wire _06387_;
  wire _06388_;
  wire _06389_;
  wire _06390_;
  wire _06391_;
  wire _06392_;
  wire _06393_;
  wire _06394_;
  wire _06395_;
  wire _06396_;
  wire _06397_;
  wire _06398_;
  wire _06399_;
  wire _06400_;
  wire _06401_;
  wire _06402_;
  wire _06403_;
  wire _06404_;
  wire _06405_;
  wire _06406_;
  wire _06407_;
  wire _06408_;
  wire _06409_;
  wire _06410_;
  wire _06411_;
  wire _06412_;
  wire _06413_;
  wire _06414_;
  wire _06415_;
  wire _06416_;
  wire _06417_;
  wire _06418_;
  wire _06419_;
  wire _06420_;
  wire _06421_;
  wire _06422_;
  wire _06423_;
  wire _06424_;
  wire _06425_;
  wire _06426_;
  wire _06427_;
  wire _06428_;
  wire _06429_;
  wire _06430_;
  wire _06431_;
  wire _06432_;
  wire _06433_;
  wire _06434_;
  wire _06435_;
  wire _06436_;
  wire _06437_;
  wire _06438_;
  wire _06439_;
  wire _06440_;
  wire _06441_;
  wire _06442_;
  wire _06443_;
  wire _06444_;
  wire _06445_;
  wire _06446_;
  wire _06447_;
  wire _06448_;
  wire _06449_;
  wire _06450_;
  wire _06451_;
  wire _06452_;
  wire _06453_;
  wire _06454_;
  wire _06455_;
  wire _06456_;
  wire _06457_;
  wire _06458_;
  wire _06459_;
  wire _06460_;
  wire _06461_;
  wire _06462_;
  wire _06463_;
  wire _06464_;
  wire _06465_;
  wire _06466_;
  wire _06467_;
  wire _06468_;
  wire _06469_;
  wire _06470_;
  wire _06471_;
  wire _06472_;
  wire _06473_;
  wire _06474_;
  wire _06475_;
  wire _06476_;
  wire _06477_;
  wire _06478_;
  wire _06479_;
  wire _06480_;
  wire _06481_;
  wire _06482_;
  wire _06483_;
  wire _06484_;
  wire _06485_;
  wire _06486_;
  wire _06487_;
  wire _06488_;
  wire _06489_;
  wire _06490_;
  wire _06491_;
  wire _06492_;
  wire _06493_;
  wire _06494_;
  wire _06495_;
  wire _06496_;
  wire _06497_;
  wire _06498_;
  wire _06499_;
  wire _06500_;
  wire _06501_;
  wire _06502_;
  wire _06503_;
  wire _06504_;
  wire _06505_;
  wire _06506_;
  wire _06507_;
  wire _06508_;
  wire _06509_;
  wire _06510_;
  wire _06511_;
  wire _06512_;
  wire _06513_;
  wire _06514_;
  wire _06515_;
  wire _06516_;
  wire _06517_;
  wire _06518_;
  wire _06519_;
  wire _06520_;
  wire _06521_;
  wire _06522_;
  wire _06523_;
  wire _06524_;
  wire _06525_;
  wire _06526_;
  wire _06527_;
  wire _06528_;
  wire _06529_;
  wire _06530_;
  wire _06531_;
  wire _06532_;
  wire _06533_;
  wire _06534_;
  wire _06535_;
  wire _06536_;
  wire _06537_;
  wire _06538_;
  wire _06539_;
  wire _06540_;
  wire _06541_;
  wire _06542_;
  wire _06543_;
  wire _06544_;
  wire _06545_;
  wire _06546_;
  wire _06547_;
  wire _06548_;
  wire _06549_;
  wire _06550_;
  wire _06551_;
  wire _06552_;
  wire _06553_;
  wire _06554_;
  wire _06555_;
  wire _06556_;
  wire _06557_;
  wire _06558_;
  wire _06559_;
  wire _06560_;
  wire _06561_;
  wire _06562_;
  wire _06563_;
  wire _06564_;
  wire _06565_;
  wire _06566_;
  wire _06567_;
  wire _06568_;
  wire _06569_;
  wire _06570_;
  wire _06571_;
  wire _06572_;
  wire _06573_;
  wire _06574_;
  wire _06575_;
  wire _06576_;
  wire _06577_;
  wire _06578_;
  wire _06579_;
  wire _06580_;
  wire _06581_;
  wire _06582_;
  wire _06583_;
  wire _06584_;
  wire _06585_;
  wire _06586_;
  wire _06587_;
  wire _06588_;
  wire _06589_;
  wire _06590_;
  wire _06591_;
  wire _06592_;
  wire _06593_;
  wire _06594_;
  wire _06595_;
  wire _06596_;
  wire _06597_;
  wire _06598_;
  wire _06599_;
  wire _06600_;
  wire _06601_;
  wire _06602_;
  wire _06603_;
  wire _06604_;
  wire _06605_;
  wire _06606_;
  wire _06607_;
  wire _06608_;
  wire _06609_;
  wire _06610_;
  wire _06611_;
  wire _06612_;
  wire _06613_;
  wire _06614_;
  wire _06615_;
  wire _06616_;
  wire _06617_;
  wire _06618_;
  wire _06619_;
  wire _06620_;
  wire _06621_;
  wire _06622_;
  wire _06623_;
  wire _06624_;
  wire _06625_;
  wire _06626_;
  wire _06627_;
  wire _06628_;
  wire _06629_;
  wire _06630_;
  wire _06631_;
  wire _06632_;
  wire _06633_;
  wire _06634_;
  wire _06635_;
  wire _06636_;
  wire _06637_;
  wire _06638_;
  wire _06639_;
  wire _06640_;
  wire _06641_;
  wire _06642_;
  wire _06643_;
  wire _06644_;
  wire _06645_;
  wire _06646_;
  wire _06647_;
  wire _06648_;
  wire _06649_;
  wire _06650_;
  wire _06651_;
  wire _06652_;
  wire _06653_;
  wire _06654_;
  wire _06655_;
  wire _06656_;
  wire _06657_;
  wire _06658_;
  wire _06659_;
  wire _06660_;
  wire _06661_;
  wire _06662_;
  wire _06663_;
  wire _06664_;
  wire _06665_;
  wire _06666_;
  wire _06667_;
  wire _06668_;
  wire _06669_;
  wire _06670_;
  wire _06671_;
  wire _06672_;
  wire _06673_;
  wire _06674_;
  wire _06675_;
  wire _06676_;
  wire _06677_;
  wire _06678_;
  wire _06679_;
  wire _06680_;
  wire _06681_;
  wire _06682_;
  wire _06683_;
  wire _06684_;
  wire _06685_;
  wire _06686_;
  wire _06687_;
  wire _06688_;
  wire _06689_;
  wire _06690_;
  wire _06691_;
  wire _06692_;
  wire _06693_;
  wire _06694_;
  wire _06695_;
  wire _06696_;
  wire _06697_;
  wire _06698_;
  wire _06699_;
  wire _06700_;
  wire _06701_;
  wire _06702_;
  wire _06703_;
  wire _06704_;
  wire _06705_;
  wire _06706_;
  wire _06707_;
  wire _06708_;
  wire _06709_;
  wire _06710_;
  wire _06711_;
  wire _06712_;
  wire _06713_;
  wire _06714_;
  wire _06715_;
  wire _06716_;
  wire _06717_;
  wire _06718_;
  wire _06719_;
  wire _06720_;
  wire _06721_;
  wire _06722_;
  wire _06723_;
  wire _06724_;
  wire _06725_;
  wire _06726_;
  wire _06727_;
  wire _06728_;
  wire _06729_;
  wire _06730_;
  wire _06731_;
  wire _06732_;
  wire _06733_;
  wire _06734_;
  wire _06735_;
  wire _06736_;
  wire _06737_;
  wire _06738_;
  wire _06739_;
  wire _06740_;
  wire _06741_;
  wire _06742_;
  wire _06743_;
  wire _06744_;
  wire _06745_;
  wire _06746_;
  wire _06747_;
  wire _06748_;
  wire _06749_;
  wire _06750_;
  wire _06751_;
  wire _06752_;
  wire _06753_;
  wire _06754_;
  wire _06755_;
  wire _06756_;
  wire _06757_;
  wire _06758_;
  wire _06759_;
  wire _06760_;
  wire _06761_;
  wire _06762_;
  wire _06763_;
  wire _06764_;
  wire _06765_;
  wire _06766_;
  wire _06767_;
  wire _06768_;
  wire _06769_;
  wire _06770_;
  wire _06771_;
  wire _06772_;
  wire _06773_;
  wire _06774_;
  wire _06775_;
  wire _06776_;
  wire _06777_;
  wire _06778_;
  wire _06779_;
  wire _06780_;
  wire _06781_;
  wire _06782_;
  wire _06783_;
  wire _06784_;
  wire _06785_;
  wire _06786_;
  wire _06787_;
  wire _06788_;
  wire _06789_;
  wire _06790_;
  wire _06791_;
  wire _06792_;
  wire _06793_;
  wire _06794_;
  wire _06795_;
  wire _06796_;
  wire _06797_;
  wire _06798_;
  wire _06799_;
  wire _06800_;
  wire _06801_;
  wire _06802_;
  wire _06803_;
  wire _06804_;
  wire _06805_;
  wire _06806_;
  wire _06807_;
  wire _06808_;
  wire _06809_;
  wire _06810_;
  wire _06811_;
  wire _06812_;
  wire _06813_;
  wire _06814_;
  wire _06815_;
  wire _06816_;
  wire _06817_;
  wire _06818_;
  wire _06819_;
  wire _06820_;
  wire _06821_;
  wire _06822_;
  wire _06823_;
  wire _06824_;
  wire _06825_;
  wire _06826_;
  wire _06827_;
  wire _06828_;
  wire _06829_;
  wire _06830_;
  wire _06831_;
  wire _06832_;
  wire _06833_;
  wire _06834_;
  wire _06835_;
  wire _06836_;
  wire _06837_;
  wire _06838_;
  wire _06839_;
  wire _06840_;
  wire _06841_;
  wire _06842_;
  wire _06843_;
  wire _06844_;
  wire _06845_;
  wire _06846_;
  wire _06847_;
  wire _06848_;
  wire _06849_;
  wire _06850_;
  wire _06851_;
  wire _06852_;
  wire _06853_;
  wire _06854_;
  wire _06855_;
  wire _06856_;
  wire _06857_;
  wire _06858_;
  wire _06859_;
  wire _06860_;
  wire _06861_;
  wire _06862_;
  wire _06863_;
  wire _06864_;
  wire _06865_;
  wire _06866_;
  wire _06867_;
  wire _06868_;
  wire _06869_;
  wire _06870_;
  wire _06871_;
  wire _06872_;
  wire _06873_;
  wire _06874_;
  wire _06875_;
  wire _06876_;
  wire _06877_;
  wire _06878_;
  wire _06879_;
  wire _06880_;
  wire _06881_;
  wire _06882_;
  wire _06883_;
  wire _06884_;
  wire _06885_;
  wire _06886_;
  wire _06887_;
  wire _06888_;
  wire _06889_;
  wire _06890_;
  wire _06891_;
  wire _06892_;
  wire _06893_;
  wire _06894_;
  wire _06895_;
  wire _06896_;
  wire _06897_;
  wire _06898_;
  wire _06899_;
  wire _06900_;
  wire _06901_;
  wire _06902_;
  wire _06903_;
  wire _06904_;
  wire _06905_;
  wire _06906_;
  wire _06907_;
  wire _06908_;
  wire _06909_;
  wire _06910_;
  wire _06911_;
  wire _06912_;
  wire _06913_;
  wire _06914_;
  wire _06915_;
  wire _06916_;
  wire _06917_;
  wire _06918_;
  wire _06919_;
  wire _06920_;
  wire _06921_;
  wire _06922_;
  wire _06923_;
  wire _06924_;
  wire _06925_;
  wire _06926_;
  wire _06927_;
  wire _06928_;
  wire _06929_;
  wire _06930_;
  wire _06931_;
  wire _06932_;
  wire _06933_;
  wire _06934_;
  wire _06935_;
  wire _06936_;
  wire _06937_;
  wire _06938_;
  wire _06939_;
  wire _06940_;
  wire _06941_;
  wire _06942_;
  wire _06943_;
  wire _06944_;
  wire _06945_;
  wire _06946_;
  wire _06947_;
  wire _06948_;
  wire _06949_;
  wire _06950_;
  wire _06951_;
  wire _06952_;
  wire _06953_;
  wire _06954_;
  wire _06955_;
  wire _06956_;
  wire _06957_;
  wire _06958_;
  wire _06959_;
  wire _06960_;
  wire _06961_;
  wire _06962_;
  wire _06963_;
  wire _06964_;
  wire _06965_;
  wire _06966_;
  wire _06967_;
  wire _06968_;
  wire _06969_;
  wire _06970_;
  wire _06971_;
  wire _06972_;
  wire _06973_;
  wire _06974_;
  wire _06975_;
  wire _06976_;
  wire _06977_;
  wire _06978_;
  wire _06979_;
  wire _06980_;
  wire _06981_;
  wire _06982_;
  wire _06983_;
  wire _06984_;
  wire _06985_;
  wire _06986_;
  wire _06987_;
  wire _06988_;
  wire _06989_;
  wire _06990_;
  wire _06991_;
  wire _06992_;
  wire _06993_;
  wire _06994_;
  wire _06995_;
  wire _06996_;
  wire _06997_;
  wire _06998_;
  wire _06999_;
  wire _07000_;
  wire _07001_;
  wire _07002_;
  wire _07003_;
  wire _07004_;
  wire _07005_;
  wire _07006_;
  wire _07007_;
  wire _07008_;
  wire _07009_;
  wire _07010_;
  wire _07011_;
  wire _07012_;
  wire _07013_;
  wire _07014_;
  wire _07015_;
  wire _07016_;
  wire _07017_;
  wire _07018_;
  wire _07019_;
  wire _07020_;
  wire _07021_;
  wire _07022_;
  wire _07023_;
  wire _07024_;
  wire _07025_;
  wire _07026_;
  wire _07027_;
  wire _07028_;
  wire _07029_;
  wire _07030_;
  wire _07031_;
  wire _07032_;
  wire _07033_;
  wire _07034_;
  wire _07035_;
  wire _07036_;
  wire _07037_;
  wire _07038_;
  wire _07039_;
  wire _07040_;
  wire _07041_;
  wire _07042_;
  wire _07043_;
  wire _07044_;
  wire _07045_;
  wire _07046_;
  wire _07047_;
  wire _07048_;
  wire _07049_;
  wire _07050_;
  wire _07051_;
  wire _07052_;
  wire _07053_;
  wire _07054_;
  wire _07055_;
  wire _07056_;
  wire _07057_;
  wire _07058_;
  wire _07059_;
  wire _07060_;
  wire _07061_;
  wire _07062_;
  wire _07063_;
  wire _07064_;
  wire _07065_;
  wire _07066_;
  wire _07067_;
  wire _07068_;
  wire _07069_;
  wire _07070_;
  wire _07071_;
  wire _07072_;
  wire _07073_;
  wire _07074_;
  wire _07075_;
  wire _07076_;
  wire _07077_;
  wire _07078_;
  wire _07079_;
  wire _07080_;
  wire _07081_;
  wire _07082_;
  wire _07083_;
  wire _07084_;
  wire _07085_;
  wire _07086_;
  wire _07087_;
  wire _07088_;
  wire _07089_;
  wire _07090_;
  wire _07091_;
  wire _07092_;
  wire _07093_;
  wire _07094_;
  wire _07095_;
  wire _07096_;
  wire _07097_;
  wire _07098_;
  wire _07099_;
  wire _07100_;
  wire _07101_;
  wire _07102_;
  wire _07103_;
  wire _07104_;
  wire _07105_;
  wire _07106_;
  wire _07107_;
  wire _07108_;
  wire _07109_;
  wire _07110_;
  wire _07111_;
  wire _07112_;
  wire _07113_;
  wire _07114_;
  wire _07115_;
  wire _07116_;
  wire _07117_;
  wire _07118_;
  wire _07119_;
  wire _07120_;
  wire _07121_;
  wire _07122_;
  wire _07123_;
  wire _07124_;
  wire _07125_;
  wire _07126_;
  wire _07127_;
  wire _07128_;
  wire _07129_;
  wire _07130_;
  wire _07131_;
  wire _07132_;
  wire _07133_;
  wire _07134_;
  wire _07135_;
  wire _07136_;
  wire _07137_;
  wire _07138_;
  wire _07139_;
  wire _07140_;
  wire _07141_;
  wire _07142_;
  wire _07143_;
  wire _07144_;
  wire _07145_;
  wire _07146_;
  wire _07147_;
  wire _07148_;
  wire _07149_;
  wire _07150_;
  wire _07151_;
  wire _07152_;
  wire _07153_;
  wire _07154_;
  wire _07155_;
  wire _07156_;
  wire _07157_;
  wire _07158_;
  wire _07159_;
  wire _07160_;
  wire _07161_;
  wire _07162_;
  wire _07163_;
  wire _07164_;
  wire _07165_;
  wire _07166_;
  wire _07167_;
  wire _07168_;
  wire _07169_;
  wire _07170_;
  wire _07171_;
  wire _07172_;
  wire _07173_;
  wire _07174_;
  wire _07175_;
  wire _07176_;
  wire _07177_;
  wire _07178_;
  wire _07179_;
  wire _07180_;
  wire _07181_;
  wire _07182_;
  wire _07183_;
  wire _07184_;
  wire _07185_;
  wire _07186_;
  wire _07187_;
  wire _07188_;
  wire _07189_;
  wire _07190_;
  wire _07191_;
  wire _07192_;
  wire _07193_;
  wire _07194_;
  wire _07195_;
  wire _07196_;
  wire _07197_;
  wire _07198_;
  wire _07199_;
  wire _07200_;
  wire _07201_;
  wire _07202_;
  wire _07203_;
  wire _07204_;
  wire _07205_;
  wire _07206_;
  wire _07207_;
  wire _07208_;
  wire _07209_;
  wire _07210_;
  wire _07211_;
  wire _07212_;
  wire _07213_;
  wire _07214_;
  wire _07215_;
  wire _07216_;
  wire _07217_;
  wire _07218_;
  wire _07219_;
  wire _07220_;
  wire _07221_;
  wire _07222_;
  wire _07223_;
  wire _07224_;
  wire _07225_;
  wire _07226_;
  wire _07227_;
  wire _07228_;
  wire _07229_;
  wire _07230_;
  wire _07231_;
  wire _07232_;
  wire _07233_;
  wire _07234_;
  wire _07235_;
  wire _07236_;
  wire _07237_;
  wire _07238_;
  wire _07239_;
  wire _07240_;
  wire _07241_;
  wire _07242_;
  wire _07243_;
  wire _07244_;
  wire _07245_;
  wire _07246_;
  wire _07247_;
  wire _07248_;
  wire _07249_;
  wire _07250_;
  wire _07251_;
  wire _07252_;
  wire _07253_;
  wire _07254_;
  wire _07255_;
  wire _07256_;
  wire _07257_;
  wire _07258_;
  wire _07259_;
  wire _07260_;
  wire _07261_;
  wire _07262_;
  wire _07263_;
  wire _07264_;
  wire _07265_;
  wire _07266_;
  wire _07267_;
  wire _07268_;
  wire _07269_;
  wire _07270_;
  wire _07271_;
  wire _07272_;
  wire _07273_;
  wire _07274_;
  wire _07275_;
  wire _07276_;
  wire _07277_;
  wire _07278_;
  wire _07279_;
  wire _07280_;
  wire _07281_;
  wire _07282_;
  wire _07283_;
  wire _07284_;
  wire _07285_;
  wire _07286_;
  wire _07287_;
  wire _07288_;
  wire _07289_;
  wire _07290_;
  wire _07291_;
  wire _07292_;
  wire _07293_;
  wire _07294_;
  wire _07295_;
  wire _07296_;
  wire _07297_;
  wire _07298_;
  wire _07299_;
  wire _07300_;
  wire _07301_;
  wire _07302_;
  wire _07303_;
  wire _07304_;
  wire _07305_;
  wire _07306_;
  wire _07307_;
  wire _07308_;
  wire _07309_;
  wire _07310_;
  wire _07311_;
  wire _07312_;
  wire _07313_;
  wire _07314_;
  wire _07315_;
  wire _07316_;
  wire _07317_;
  wire _07318_;
  wire _07319_;
  wire _07320_;
  wire _07321_;
  wire _07322_;
  wire _07323_;
  wire _07324_;
  wire _07325_;
  wire _07326_;
  wire _07327_;
  wire _07328_;
  wire _07329_;
  wire _07330_;
  wire _07331_;
  wire _07332_;
  wire _07333_;
  wire _07334_;
  wire _07335_;
  wire _07336_;
  wire _07337_;
  wire _07338_;
  wire _07339_;
  wire _07340_;
  wire _07341_;
  wire _07342_;
  wire _07343_;
  wire _07344_;
  wire _07345_;
  wire _07346_;
  wire _07347_;
  wire _07348_;
  wire _07349_;
  wire _07350_;
  wire _07351_;
  wire _07352_;
  wire _07353_;
  wire _07354_;
  wire _07355_;
  wire _07356_;
  wire _07357_;
  wire _07358_;
  wire _07359_;
  wire _07360_;
  wire _07361_;
  wire _07362_;
  wire _07363_;
  wire _07364_;
  wire _07365_;
  wire _07366_;
  wire _07367_;
  wire _07368_;
  wire _07369_;
  wire _07370_;
  wire _07371_;
  wire _07372_;
  wire _07373_;
  wire _07374_;
  wire _07375_;
  wire _07376_;
  wire _07377_;
  wire _07378_;
  wire _07379_;
  wire _07380_;
  wire _07381_;
  wire _07382_;
  wire _07383_;
  wire _07384_;
  wire _07385_;
  wire _07386_;
  wire _07387_;
  wire _07388_;
  wire _07389_;
  wire _07390_;
  wire _07391_;
  wire _07392_;
  wire _07393_;
  wire _07394_;
  wire _07395_;
  wire _07396_;
  wire _07397_;
  wire _07398_;
  wire _07399_;
  wire _07400_;
  wire _07401_;
  wire _07402_;
  wire _07403_;
  wire _07404_;
  wire _07405_;
  wire _07406_;
  wire _07407_;
  wire _07408_;
  wire _07409_;
  wire _07410_;
  wire _07411_;
  wire _07412_;
  wire _07413_;
  wire _07414_;
  wire _07415_;
  wire _07416_;
  wire _07417_;
  wire _07418_;
  wire _07419_;
  wire _07420_;
  wire _07421_;
  wire _07422_;
  wire _07423_;
  wire _07424_;
  wire _07425_;
  wire _07426_;
  wire _07427_;
  wire _07428_;
  wire _07429_;
  wire _07430_;
  wire _07431_;
  wire _07432_;
  wire _07433_;
  wire _07434_;
  wire _07435_;
  wire _07436_;
  wire _07437_;
  wire _07438_;
  wire _07439_;
  wire _07440_;
  wire _07441_;
  wire _07442_;
  wire _07443_;
  wire _07444_;
  wire _07445_;
  wire _07446_;
  wire _07447_;
  wire _07448_;
  wire _07449_;
  wire _07450_;
  wire _07451_;
  wire _07452_;
  wire _07453_;
  wire _07454_;
  wire _07455_;
  wire _07456_;
  wire _07457_;
  wire _07458_;
  wire _07459_;
  wire _07460_;
  wire _07461_;
  wire _07462_;
  wire _07463_;
  wire _07464_;
  wire _07465_;
  wire _07466_;
  wire _07467_;
  wire _07468_;
  wire _07469_;
  wire _07470_;
  wire _07471_;
  wire _07472_;
  wire _07473_;
  wire _07474_;
  wire _07475_;
  wire _07476_;
  wire _07477_;
  wire _07478_;
  wire _07479_;
  wire _07480_;
  wire _07481_;
  wire _07482_;
  wire _07483_;
  wire _07484_;
  wire _07485_;
  wire _07486_;
  wire _07487_;
  wire _07488_;
  wire _07489_;
  wire _07490_;
  wire _07491_;
  wire _07492_;
  wire _07493_;
  wire _07494_;
  wire _07495_;
  wire _07496_;
  wire _07497_;
  wire _07498_;
  wire _07499_;
  wire _07500_;
  wire _07501_;
  wire _07502_;
  wire _07503_;
  wire _07504_;
  wire _07505_;
  wire _07506_;
  wire _07507_;
  wire _07508_;
  wire _07509_;
  wire _07510_;
  wire _07511_;
  wire _07512_;
  wire _07513_;
  wire _07514_;
  wire _07515_;
  wire _07516_;
  wire _07517_;
  wire _07518_;
  wire _07519_;
  wire _07520_;
  wire _07521_;
  wire _07522_;
  wire _07523_;
  wire _07524_;
  wire _07525_;
  wire _07526_;
  wire _07527_;
  wire _07528_;
  wire _07529_;
  wire _07530_;
  wire _07531_;
  wire _07532_;
  wire _07533_;
  wire _07534_;
  wire _07535_;
  wire _07536_;
  wire _07537_;
  wire _07538_;
  wire _07539_;
  wire _07540_;
  wire _07541_;
  wire _07542_;
  wire _07543_;
  wire _07544_;
  wire _07545_;
  wire _07546_;
  wire _07547_;
  wire _07548_;
  wire _07549_;
  wire _07550_;
  wire _07551_;
  wire _07552_;
  wire _07553_;
  wire _07554_;
  wire _07555_;
  wire _07556_;
  wire _07557_;
  wire _07558_;
  wire _07559_;
  wire _07560_;
  wire _07561_;
  wire _07562_;
  wire _07563_;
  wire _07564_;
  wire _07565_;
  wire _07566_;
  wire _07567_;
  wire _07568_;
  wire _07569_;
  wire _07570_;
  wire _07571_;
  wire _07572_;
  wire _07573_;
  wire _07574_;
  wire _07575_;
  wire _07576_;
  wire _07577_;
  wire _07578_;
  wire _07579_;
  wire _07580_;
  wire _07581_;
  wire _07582_;
  wire _07583_;
  wire _07584_;
  wire _07585_;
  wire _07586_;
  wire _07587_;
  wire _07588_;
  wire _07589_;
  wire _07590_;
  wire _07591_;
  wire _07592_;
  wire _07593_;
  wire _07594_;
  wire _07595_;
  wire _07596_;
  wire _07597_;
  wire _07598_;
  wire _07599_;
  wire _07600_;
  wire _07601_;
  wire _07602_;
  wire _07603_;
  wire _07604_;
  wire _07605_;
  wire _07606_;
  wire _07607_;
  wire _07608_;
  wire _07609_;
  wire _07610_;
  wire _07611_;
  wire _07612_;
  wire _07613_;
  wire _07614_;
  wire _07615_;
  wire _07616_;
  wire _07617_;
  wire _07618_;
  wire _07619_;
  wire _07620_;
  wire _07621_;
  wire _07622_;
  wire _07623_;
  wire _07624_;
  wire _07625_;
  wire _07626_;
  wire _07627_;
  wire _07628_;
  wire _07629_;
  wire _07630_;
  wire _07631_;
  wire _07632_;
  wire _07633_;
  wire _07634_;
  wire _07635_;
  wire _07636_;
  wire _07637_;
  wire _07638_;
  wire _07639_;
  wire _07640_;
  wire _07641_;
  wire _07642_;
  wire _07643_;
  wire _07644_;
  wire _07645_;
  wire _07646_;
  wire _07647_;
  wire _07648_;
  wire _07649_;
  wire _07650_;
  wire _07651_;
  wire _07652_;
  wire _07653_;
  wire _07654_;
  wire _07655_;
  wire _07656_;
  wire _07657_;
  wire _07658_;
  wire _07659_;
  wire _07660_;
  wire _07661_;
  wire _07662_;
  wire _07663_;
  wire _07664_;
  wire _07665_;
  wire _07666_;
  wire _07667_;
  wire _07668_;
  wire _07669_;
  wire _07670_;
  wire _07671_;
  wire _07672_;
  wire _07673_;
  wire _07674_;
  wire _07675_;
  wire _07676_;
  wire _07677_;
  wire _07678_;
  wire _07679_;
  wire _07680_;
  wire _07681_;
  wire _07682_;
  wire _07683_;
  wire _07684_;
  wire _07685_;
  wire _07686_;
  wire _07687_;
  wire _07688_;
  wire _07689_;
  wire _07690_;
  wire _07691_;
  wire _07692_;
  wire _07693_;
  wire _07694_;
  wire _07695_;
  wire _07696_;
  wire _07697_;
  wire _07698_;
  wire _07699_;
  wire _07700_;
  wire _07701_;
  wire _07702_;
  wire _07703_;
  wire _07704_;
  wire _07705_;
  wire _07706_;
  wire _07707_;
  wire _07708_;
  wire _07709_;
  wire _07710_;
  wire _07711_;
  wire _07712_;
  wire _07713_;
  wire _07714_;
  wire _07715_;
  wire _07716_;
  wire _07717_;
  wire _07718_;
  wire _07719_;
  wire _07720_;
  wire _07721_;
  wire _07722_;
  wire _07723_;
  wire _07724_;
  wire _07725_;
  wire _07726_;
  wire _07727_;
  wire _07728_;
  wire _07729_;
  wire _07730_;
  wire _07731_;
  wire _07732_;
  wire _07733_;
  wire _07734_;
  wire _07735_;
  wire _07736_;
  wire _07737_;
  wire _07738_;
  wire _07739_;
  wire _07740_;
  wire _07741_;
  wire _07742_;
  wire _07743_;
  wire _07744_;
  wire _07745_;
  wire _07746_;
  wire _07747_;
  wire _07748_;
  wire _07749_;
  wire _07750_;
  wire _07751_;
  wire _07752_;
  wire _07753_;
  wire _07754_;
  wire _07755_;
  wire _07756_;
  wire _07757_;
  wire _07758_;
  wire _07759_;
  wire _07760_;
  wire _07761_;
  wire _07762_;
  wire _07763_;
  wire _07764_;
  wire _07765_;
  wire _07766_;
  wire _07767_;
  wire _07768_;
  wire _07769_;
  wire _07770_;
  wire _07771_;
  wire _07772_;
  wire _07773_;
  wire _07774_;
  wire _07775_;
  wire _07776_;
  wire _07777_;
  wire _07778_;
  wire _07779_;
  wire _07780_;
  wire _07781_;
  wire _07782_;
  wire _07783_;
  wire _07784_;
  wire _07785_;
  wire _07786_;
  wire _07787_;
  wire _07788_;
  wire _07789_;
  wire _07790_;
  wire _07791_;
  wire _07792_;
  wire _07793_;
  wire _07794_;
  wire _07795_;
  wire _07796_;
  wire _07797_;
  wire _07798_;
  wire _07799_;
  wire _07800_;
  wire _07801_;
  wire _07802_;
  wire _07803_;
  wire _07804_;
  wire _07805_;
  wire _07806_;
  wire _07807_;
  wire _07808_;
  wire _07809_;
  wire _07810_;
  wire _07811_;
  wire _07812_;
  wire _07813_;
  wire _07814_;
  wire _07815_;
  wire _07816_;
  wire _07817_;
  wire _07818_;
  wire _07819_;
  wire _07820_;
  wire _07821_;
  wire _07822_;
  wire _07823_;
  wire _07824_;
  wire _07825_;
  wire _07826_;
  wire _07827_;
  wire _07828_;
  wire _07829_;
  wire _07830_;
  wire _07831_;
  wire _07832_;
  wire _07833_;
  wire _07834_;
  wire _07835_;
  wire _07836_;
  wire _07837_;
  wire _07838_;
  wire _07839_;
  wire _07840_;
  wire _07841_;
  wire _07842_;
  wire _07843_;
  wire _07844_;
  wire _07845_;
  wire _07846_;
  wire _07847_;
  wire _07848_;
  wire _07849_;
  wire _07850_;
  wire _07851_;
  wire _07852_;
  wire _07853_;
  wire _07854_;
  wire _07855_;
  wire _07856_;
  wire _07857_;
  wire _07858_;
  wire _07859_;
  wire _07860_;
  wire _07861_;
  wire _07862_;
  wire _07863_;
  wire _07864_;
  wire _07865_;
  wire _07866_;
  wire _07867_;
  wire _07868_;
  wire _07869_;
  wire _07870_;
  wire _07871_;
  wire _07872_;
  wire _07873_;
  wire _07874_;
  wire _07875_;
  wire _07876_;
  wire _07877_;
  wire _07878_;
  wire _07879_;
  wire _07880_;
  wire _07881_;
  wire _07882_;
  wire _07883_;
  wire _07884_;
  wire _07885_;
  wire _07886_;
  wire _07887_;
  wire _07888_;
  wire _07889_;
  wire _07890_;
  wire _07891_;
  wire _07892_;
  wire _07893_;
  wire _07894_;
  wire _07895_;
  wire _07896_;
  wire _07897_;
  wire _07898_;
  wire _07899_;
  wire _07900_;
  wire _07901_;
  wire _07902_;
  wire _07903_;
  wire _07904_;
  wire _07905_;
  wire _07906_;
  wire _07907_;
  wire _07908_;
  wire _07909_;
  wire _07910_;
  wire _07911_;
  wire _07912_;
  wire _07913_;
  wire _07914_;
  wire _07915_;
  wire _07916_;
  wire _07917_;
  wire _07918_;
  wire _07919_;
  wire _07920_;
  wire _07921_;
  wire _07922_;
  wire _07923_;
  wire _07924_;
  wire _07925_;
  wire _07926_;
  wire _07927_;
  wire _07928_;
  wire _07929_;
  wire _07930_;
  wire _07931_;
  wire _07932_;
  wire _07933_;
  wire _07934_;
  wire _07935_;
  wire _07936_;
  wire _07937_;
  wire _07938_;
  wire _07939_;
  wire _07940_;
  wire _07941_;
  wire _07942_;
  wire _07943_;
  wire _07944_;
  wire _07945_;
  wire _07946_;
  wire _07947_;
  wire _07948_;
  wire _07949_;
  wire _07950_;
  wire _07951_;
  wire _07952_;
  wire _07953_;
  wire _07954_;
  wire _07955_;
  wire _07956_;
  wire _07957_;
  wire _07958_;
  wire _07959_;
  wire _07960_;
  wire _07961_;
  wire _07962_;
  wire _07963_;
  wire _07964_;
  wire _07965_;
  wire _07966_;
  wire _07967_;
  wire _07968_;
  wire _07969_;
  wire _07970_;
  wire _07971_;
  wire _07972_;
  wire _07973_;
  wire _07974_;
  wire _07975_;
  wire _07976_;
  wire _07977_;
  wire _07978_;
  wire _07979_;
  wire _07980_;
  wire _07981_;
  wire _07982_;
  wire _07983_;
  wire _07984_;
  wire _07985_;
  wire _07986_;
  wire _07987_;
  wire _07988_;
  wire _07989_;
  wire _07990_;
  wire _07991_;
  wire _07992_;
  wire _07993_;
  wire _07994_;
  wire _07995_;
  wire _07996_;
  wire _07997_;
  wire _07998_;
  wire _07999_;
  wire _08000_;
  input MemRead_i;
  input MemWrite_i;
  input \addr_i[0];
  input \addr_i[10];
  input \addr_i[11];
  input \addr_i[12];
  input \addr_i[13];
  input \addr_i[14];
  input \addr_i[15];
  input \addr_i[16];
  input \addr_i[17];
  input \addr_i[18];
  input \addr_i[19];
  input \addr_i[1];
  input \addr_i[20];
  input \addr_i[21];
  input \addr_i[22];
  input \addr_i[23];
  input \addr_i[24];
  input \addr_i[25];
  input \addr_i[26];
  input \addr_i[27];
  input \addr_i[28];
  input \addr_i[29];
  input \addr_i[2];
  input \addr_i[30];
  input \addr_i[31];
  input \addr_i[3];
  input \addr_i[4];
  input \addr_i[5];
  input \addr_i[6];
  input \addr_i[7];
  input \addr_i[8];
  input \addr_i[9];
  input \data_i[0];
  input \data_i[10];
  input \data_i[11];
  input \data_i[12];
  input \data_i[13];
  input \data_i[14];
  input \data_i[15];
  input \data_i[16];
  input \data_i[17];
  input \data_i[18];
  input \data_i[19];
  input \data_i[1];
  input \data_i[20];
  input \data_i[21];
  input \data_i[22];
  input \data_i[23];
  input \data_i[24];
  input \data_i[25];
  input \data_i[26];
  input \data_i[27];
  input \data_i[28];
  input \data_i[29];
  input \data_i[2];
  input \data_i[30];
  input \data_i[31];
  input \data_i[3];
  input \data_i[4];
  input \data_i[5];
  input \data_i[6];
  input \data_i[7];
  input \data_i[8];
  input \data_i[9];
  input \memory[0][0];
  input \memory[0][1];
  input \memory[0][2];
  input \memory[0][3];
  input \memory[0][4];
  input \memory[0][5];
  input \memory[0][6];
  input \memory[0][7];
  input \memory[10][0];
  input \memory[10][1];
  input \memory[10][2];
  input \memory[10][3];
  input \memory[10][4];
  input \memory[10][5];
  input \memory[10][6];
  input \memory[10][7];
  input \memory[11][0];
  input \memory[11][1];
  input \memory[11][2];
  input \memory[11][3];
  input \memory[11][4];
  input \memory[11][5];
  input \memory[11][6];
  input \memory[11][7];
  input \memory[12][0];
  input \memory[12][1];
  input \memory[12][2];
  input \memory[12][3];
  input \memory[12][4];
  input \memory[12][5];
  input \memory[12][6];
  input \memory[12][7];
  input \memory[13][0];
  input \memory[13][1];
  input \memory[13][2];
  input \memory[13][3];
  input \memory[13][4];
  input \memory[13][5];
  input \memory[13][6];
  input \memory[13][7];
  input \memory[14][0];
  input \memory[14][1];
  input \memory[14][2];
  input \memory[14][3];
  input \memory[14][4];
  input \memory[14][5];
  input \memory[14][6];
  input \memory[14][7];
  input \memory[15][0];
  input \memory[15][1];
  input \memory[15][2];
  input \memory[15][3];
  input \memory[15][4];
  input \memory[15][5];
  input \memory[15][6];
  input \memory[15][7];
  input \memory[16][0];
  input \memory[16][1];
  input \memory[16][2];
  input \memory[16][3];
  input \memory[16][4];
  input \memory[16][5];
  input \memory[16][6];
  input \memory[16][7];
  input \memory[17][0];
  input \memory[17][1];
  input \memory[17][2];
  input \memory[17][3];
  input \memory[17][4];
  input \memory[17][5];
  input \memory[17][6];
  input \memory[17][7];
  input \memory[18][0];
  input \memory[18][1];
  input \memory[18][2];
  input \memory[18][3];
  input \memory[18][4];
  input \memory[18][5];
  input \memory[18][6];
  input \memory[18][7];
  input \memory[19][0];
  input \memory[19][1];
  input \memory[19][2];
  input \memory[19][3];
  input \memory[19][4];
  input \memory[19][5];
  input \memory[19][6];
  input \memory[19][7];
  input \memory[1][0];
  input \memory[1][1];
  input \memory[1][2];
  input \memory[1][3];
  input \memory[1][4];
  input \memory[1][5];
  input \memory[1][6];
  input \memory[1][7];
  input \memory[20][0];
  input \memory[20][1];
  input \memory[20][2];
  input \memory[20][3];
  input \memory[20][4];
  input \memory[20][5];
  input \memory[20][6];
  input \memory[20][7];
  input \memory[21][0];
  input \memory[21][1];
  input \memory[21][2];
  input \memory[21][3];
  input \memory[21][4];
  input \memory[21][5];
  input \memory[21][6];
  input \memory[21][7];
  input \memory[22][0];
  input \memory[22][1];
  input \memory[22][2];
  input \memory[22][3];
  input \memory[22][4];
  input \memory[22][5];
  input \memory[22][6];
  input \memory[22][7];
  input \memory[23][0];
  input \memory[23][1];
  input \memory[23][2];
  input \memory[23][3];
  input \memory[23][4];
  input \memory[23][5];
  input \memory[23][6];
  input \memory[23][7];
  input \memory[24][0];
  input \memory[24][1];
  input \memory[24][2];
  input \memory[24][3];
  input \memory[24][4];
  input \memory[24][5];
  input \memory[24][6];
  input \memory[24][7];
  input \memory[25][0];
  input \memory[25][1];
  input \memory[25][2];
  input \memory[25][3];
  input \memory[25][4];
  input \memory[25][5];
  input \memory[25][6];
  input \memory[25][7];
  input \memory[26][0];
  input \memory[26][1];
  input \memory[26][2];
  input \memory[26][3];
  input \memory[26][4];
  input \memory[26][5];
  input \memory[26][6];
  input \memory[26][7];
  input \memory[27][0];
  input \memory[27][1];
  input \memory[27][2];
  input \memory[27][3];
  input \memory[27][4];
  input \memory[27][5];
  input \memory[27][6];
  input \memory[27][7];
  input \memory[28][0];
  input \memory[28][1];
  input \memory[28][2];
  input \memory[28][3];
  input \memory[28][4];
  input \memory[28][5];
  input \memory[28][6];
  input \memory[28][7];
  input \memory[29][0];
  input \memory[29][1];
  input \memory[29][2];
  input \memory[29][3];
  input \memory[29][4];
  input \memory[29][5];
  input \memory[29][6];
  input \memory[29][7];
  input \memory[2][0];
  input \memory[2][1];
  input \memory[2][2];
  input \memory[2][3];
  input \memory[2][4];
  input \memory[2][5];
  input \memory[2][6];
  input \memory[2][7];
  input \memory[30][0];
  input \memory[30][1];
  input \memory[30][2];
  input \memory[30][3];
  input \memory[30][4];
  input \memory[30][5];
  input \memory[30][6];
  input \memory[30][7];
  input \memory[31][0];
  input \memory[31][1];
  input \memory[31][2];
  input \memory[31][3];
  input \memory[31][4];
  input \memory[31][5];
  input \memory[31][6];
  input \memory[31][7];
  input \memory[3][0];
  input \memory[3][1];
  input \memory[3][2];
  input \memory[3][3];
  input \memory[3][4];
  input \memory[3][5];
  input \memory[3][6];
  input \memory[3][7];
  input \memory[4][0];
  input \memory[4][1];
  input \memory[4][2];
  input \memory[4][3];
  input \memory[4][4];
  input \memory[4][5];
  input \memory[4][6];
  input \memory[4][7];
  input \memory[5][0];
  input \memory[5][1];
  input \memory[5][2];
  input \memory[5][3];
  input \memory[5][4];
  input \memory[5][5];
  input \memory[5][6];
  input \memory[5][7];
  input \memory[6][0];
  input \memory[6][1];
  input \memory[6][2];
  input \memory[6][3];
  input \memory[6][4];
  input \memory[6][5];
  input \memory[6][6];
  input \memory[6][7];
  input \memory[7][0];
  input \memory[7][1];
  input \memory[7][2];
  input \memory[7][3];
  input \memory[7][4];
  input \memory[7][5];
  input \memory[7][6];
  input \memory[7][7];
  input \memory[8][0];
  input \memory[8][1];
  input \memory[8][2];
  input \memory[8][3];
  input \memory[8][4];
  input \memory[8][5];
  input \memory[8][6];
  input \memory[8][7];
  input \memory[9][0];
  input \memory[9][1];
  input \memory[9][2];
  input \memory[9][3];
  input \memory[9][4];
  input \memory[9][5];
  input \memory[9][6];
  input \memory[9][7];
  input \op_addr[0];
  input \op_addr[1];
  input \op_addr[2];
  input \op_addr[3];
  input \op_addr[4];
  input clk_i;
  input reset;
  output \data_mem_o[0];
  output \data_mem_o[10];
  output \data_mem_o[11];
  output \data_mem_o[12];
  output \data_mem_o[13];
  output \data_mem_o[14];
  output \data_mem_o[15];
  output \data_mem_o[16];
  output \data_mem_o[17];
  output \data_mem_o[18];
  output \data_mem_o[19];
  output \data_mem_o[1];
  output \data_mem_o[20];
  output \data_mem_o[21];
  output \data_mem_o[22];
  output \data_mem_o[23];
  output \data_mem_o[24];
  output \data_mem_o[25];
  output \data_mem_o[26];
  output \data_mem_o[27];
  output \data_mem_o[28];
  output \data_mem_o[29];
  output \data_mem_o[2];
  output \data_mem_o[30];
  output \data_mem_o[31];
  output \data_mem_o[3];
  output \data_mem_o[4];
  output \data_mem_o[5];
  output \data_mem_o[6];
  output \data_mem_o[7];
  output \data_mem_o[8];
  output \data_mem_o[9];
  output \data_o[0];
  output \data_o[10];
  output \data_o[11];
  output \data_o[12];
  output \data_o[13];
  output \data_o[14];
  output \data_o[15];
  output \data_o[16];
  output \data_o[17];
  output \data_o[18];
  output \data_o[19];
  output \data_o[1];
  output \data_o[20];
  output \data_o[21];
  output \data_o[22];
  output \data_o[23];
  output \data_o[24];
  output \data_o[25];
  output \data_o[26];
  output \data_o[27];
  output \data_o[28];
  output \data_o[29];
  output \data_o[2];
  output \data_o[30];
  output \data_o[31];
  output \data_o[3];
  output \data_o[4];
  output \data_o[5];
  output \data_o[6];
  output \data_o[7];
  output \data_o[8];
  output \data_o[9];
  output _00000_;
  output _00001_;
  output _00002_;
  output _00003_;
  output _00004_;
  output _00005_;
  output _00006_;
  output _00007_;
  output _00008_;
  output _00009_;
  output _00010_;
  output _00011_;
  output _00012_;
  output _00013_;
  output _00014_;
  output _00015_;
  output _00016_;
  output _00017_;
  output _00018_;
  output _00019_;
  output _00020_;
  output _00021_;
  output _00022_;
  output _00023_;
  output _00024_;
  output _00025_;
  output _00026_;
  output _00027_;
  output _00028_;
  output _00029_;
  output _00030_;
  output _00031_;
  output _00032_;
  output _00033_;
  output _00034_;
  output _00035_;
  output _00036_;
  output _00037_;
  output _00038_;
  output _00039_;
  output _00040_;
  output _00041_;
  output _00042_;
  output _00043_;
  output _00044_;
  output _00045_;
  output _00046_;
  output _00047_;
  output _00048_;
  output _00049_;
  output _00050_;
  output _00051_;
  output _00052_;
  output _00053_;
  output _00054_;
  output _00055_;
  output _00056_;
  output _00057_;
  output _00058_;
  output _00059_;
  output _00060_;
  output _00061_;
  output _00062_;
  output _00063_;
  output _00064_;
  output _00065_;
  output _00066_;
  output _00067_;
  output _00068_;
  output _00069_;
  output _00070_;
  output _00071_;
  output _00072_;
  output _00073_;
  output _00074_;
  output _00075_;
  output _00076_;
  output _00077_;
  output _00078_;
  output _00079_;
  output _00080_;
  output _00081_;
  output _00082_;
  output _00083_;
  output _00084_;
  output _00085_;
  output _00086_;
  output _00087_;
  output _00088_;
  output _00089_;
  output _00090_;
  output _00091_;
  output _00092_;
  output _00093_;
  output _00094_;
  output _00095_;
  output _00096_;
  output _00097_;
  output _00098_;
  output _00099_;
  output _00100_;
  output _00101_;
  output _00102_;
  output _00103_;
  output _00104_;
  output _00105_;
  output _00106_;
  output _00107_;
  output _00108_;
  output _00109_;
  output _00110_;
  output _00111_;
  output _00112_;
  output _00113_;
  output _00114_;
  output _00115_;
  output _00116_;
  output _00117_;
  output _00118_;
  output _00119_;
  output _00120_;
  output _00121_;
  output _00122_;
  output _00123_;
  output _00124_;
  output _00125_;
  output _00126_;
  output _00127_;
  output _00128_;
  output _00129_;
  output _00130_;
  output _00131_;
  output _00132_;
  output _00133_;
  output _00134_;
  output _00135_;
  output _00136_;
  output _00137_;
  output _00138_;
  output _00139_;
  output _00140_;
  output _00141_;
  output _00142_;
  output _00143_;
  output _00144_;
  output _00145_;
  output _00146_;
  output _00147_;
  output _00148_;
  output _00149_;
  output _00150_;
  output _00151_;
  output _00152_;
  output _00153_;
  output _00154_;
  output _00155_;
  output _00156_;
  output _00157_;
  output _00158_;
  output _00159_;
  output _00160_;
  output _00161_;
  output _00162_;
  output _00163_;
  output _00164_;
  output _00165_;
  output _00166_;
  output _00167_;
  output _00168_;
  output _00169_;
  output _00170_;
  output _00171_;
  output _00172_;
  output _00173_;
  output _00174_;
  output _00175_;
  output _00176_;
  output _00177_;
  output _00178_;
  output _00179_;
  output _00180_;
  output _00181_;
  output _00182_;
  output _00183_;
  output _00184_;
  output _00185_;
  output _00186_;
  output _00187_;
  output _00188_;
  output _00189_;
  output _00190_;
  output _00191_;
  output _00192_;
  output _00193_;
  output _00194_;
  output _00195_;
  output _00196_;
  output _00197_;
  output _00198_;
  output _00199_;
  output _00200_;
  output _00201_;
  output _00202_;
  output _00203_;
  output _00204_;
  output _00205_;
  output _00206_;
  output _00207_;
  output _00208_;
  output _00209_;
  output _00210_;
  output _00211_;
  output _00212_;
  output _00213_;
  output _00214_;
  output _00215_;
  output _00216_;
  output _00217_;
  output _00218_;
  output _00219_;
  output _00220_;
  output _00221_;
  output _00222_;
  output _00223_;
  output _00224_;
  output _00225_;
  output _00226_;
  output _00227_;
  output _00228_;
  output _00229_;
  output _00230_;
  output _00231_;
  output _00232_;
  output _00233_;
  output _00234_;
  output _00235_;
  output _00236_;
  output _00237_;
  output _00238_;
  output _00239_;
  output _00240_;
  output _00241_;
  output _00242_;
  output _00243_;
  output _00244_;
  output _00245_;
  output _00246_;
  output _00247_;
  output _00248_;
  output _00249_;
  output _00250_;
  output _00251_;
  output _00252_;
  output _00253_;
  output _00254_;
  output _00255_;
  AND _08008_ (
    .A(\op_addr[1] ),
    .B(\op_addr[2] ),
    .Y(_05372_)
  );
  AND _08009_ (
    .A(\op_addr[3] ),
    .B(_05372_),
    .Y(_05382_)
  );
  AND _08010_ (
    .A(_05310_),
    .B(_05382_),
    .Y(_05392_)
  );
  XOR _08011_ (
    .A(\op_addr[4] ),
    .B(_05382_),
    .Y(_05403_)
  );
  XOR _08012_ (
    .A(\op_addr[1] ),
    .B(\op_addr[2] ),
    .Y(_05413_)
  );
  AND _08014_ (
    .A(_05299_),
    .B(_05413_),
    .Y(_05434_)
  );
  NOR _08015_ (
    .A(\op_addr[1] ),
    .B(_05320_),
    .Y(_05444_)
  );
  AND _08016_ (
    .A(_05434_),
    .B(_05444_),
    .Y(_05454_)
  );
  NAND _08017_ (
    .A(_05434_),
    .B(_05444_),
    .Y(_05465_)
  );
  NOR _08018_ (
    .A(_05403_),
    .B(_05465_),
    .Y(_05475_)
  );
  NAND _08019_ (
    .A(\memory[7][0] ),
    .B(_05475_),
    .Y(_05485_)
  );
  NOR _08020_ (
    .A(\op_addr[1] ),
    .B(\op_addr[0] ),
    .Y(_05496_)
  );
  NOR _08021_ (
    .A(\op_addr[2] ),
    .B(\op_addr[3] ),
    .Y(_05506_)
  );
  XOR _08022_ (
    .A(\op_addr[3] ),
    .B(_05372_),
    .Y(_05516_)
  );
  NOR _08023_ (
    .A(_05413_),
    .B(_05516_),
    .Y(_05527_)
  );
  AND _08024_ (
    .A(_05496_),
    .B(_05506_),
    .Y(_05537_)
  );
  NAND _08025_ (
    .A(_05496_),
    .B(_05506_),
    .Y(_05547_)
  );
  AND _08026_ (
    .A(_05403_),
    .B(_05537_),
    .Y(_05558_)
  );
  NAND _08027_ (
    .A(\memory[18][0] ),
    .B(_05558_),
    .Y(_05568_)
  );
  AND _08028_ (
    .A(_05444_),
    .B(_05506_),
    .Y(_05578_)
  );
  NAND _08029_ (
    .A(_05444_),
    .B(_05506_),
    .Y(_05589_)
  );
  NOR _08030_ (
    .A(_05403_),
    .B(_05589_),
    .Y(_05599_)
  );
  NAND _08031_ (
    .A(\memory[3][0] ),
    .B(_05599_),
    .Y(_05609_)
  );
  AND _08032_ (
    .A(\op_addr[1] ),
    .B(_05320_),
    .Y(_05620_)
  );
  AND _08034_ (
    .A(\op_addr[3] ),
    .B(_05413_),
    .Y(_05640_)
  );
  AND _08035_ (
    .A(_05310_),
    .B(_05640_),
    .Y(_05651_)
  );
  AND _08036_ (
    .A(_05620_),
    .B(_05651_),
    .Y(_05661_)
  );
  NAND _08037_ (
    .A(\memory[12][0] ),
    .B(_05661_),
    .Y(_05671_)
  );
  AND _08038_ (
    .A(\op_addr[4] ),
    .B(_05640_),
    .Y(_05682_)
  );
  AND _08039_ (
    .A(_05444_),
    .B(_05682_),
    .Y(_05692_)
  );
  NAND _08040_ (
    .A(\memory[31][0] ),
    .B(_05692_),
    .Y(_05702_)
  );
  AND _08041_ (
    .A(_05434_),
    .B(_05496_),
    .Y(_05713_)
  );
  NAND _08042_ (
    .A(_05434_),
    .B(_05496_),
    .Y(_05723_)
  );
  NOR _08043_ (
    .A(_05403_),
    .B(_05723_),
    .Y(_05733_)
  );
  NAND _08044_ (
    .A(\memory[6][0] ),
    .B(_05733_),
    .Y(_05744_)
  );
  AND _08045_ (
    .A(_05403_),
    .B(_05578_),
    .Y(_05754_)
  );
  NAND _08046_ (
    .A(\memory[19][0] ),
    .B(_05754_),
    .Y(_05764_)
  );
  AND _08047_ (
    .A(\op_addr[1] ),
    .B(\op_addr[0] ),
    .Y(_05775_)
  );
  AND _08048_ (
    .A(_05651_),
    .B(_05775_),
    .Y(_05785_)
  );
  NAND _08049_ (
    .A(\memory[13][0] ),
    .B(_05785_),
    .Y(_05795_)
  );
  AND _08050_ (
    .A(_05403_),
    .B(_05713_),
    .Y(_05806_)
  );
  NAND _08051_ (
    .A(\memory[22][0] ),
    .B(_05806_),
    .Y(_05816_)
  );
  AND _08052_ (
    .A(_05496_),
    .B(_05682_),
    .Y(_05826_)
  );
  NAND _08053_ (
    .A(\memory[30][0] ),
    .B(_05826_),
    .Y(_05837_)
  );
  AND _08054_ (
    .A(_05682_),
    .B(_05775_),
    .Y(_05847_)
  );
  NAND _08055_ (
    .A(\memory[29][0] ),
    .B(_05847_),
    .Y(_05857_)
  );
  AND _08056_ (
    .A(_05423_),
    .B(_05516_),
    .Y(_05868_)
  );
  AND _08057_ (
    .A(_05496_),
    .B(_05868_),
    .Y(_05878_)
  );
  NAND _08058_ (
    .A(_05496_),
    .B(_05868_),
    .Y(_05888_)
  );
  NOR _08059_ (
    .A(_05403_),
    .B(_05888_),
    .Y(_05899_)
  );
  NAND _08060_ (
    .A(\memory[10][0] ),
    .B(_05899_),
    .Y(_05909_)
  );
  AND _08061_ (
    .A(_05403_),
    .B(_05620_),
    .Y(_05919_)
  );
  AND _08062_ (
    .A(_05434_),
    .B(_05919_),
    .Y(_05930_)
  );
  NAND _08063_ (
    .A(\memory[20][0] ),
    .B(_05930_),
    .Y(_05940_)
  );
  NOR _08064_ (
    .A(_05403_),
    .B(_05630_),
    .Y(_05950_)
  );
  AND _08065_ (
    .A(_05434_),
    .B(_05950_),
    .Y(_05961_)
  );
  NAND _08066_ (
    .A(\memory[4][0] ),
    .B(_05961_),
    .Y(_05971_)
  );
  AND _08067_ (
    .A(_05640_),
    .B(_05919_),
    .Y(_05981_)
  );
  NAND _08068_ (
    .A(\memory[28][0] ),
    .B(_05981_),
    .Y(_05992_)
  );
  AND _08069_ (
    .A(_05496_),
    .B(_05651_),
    .Y(_06002_)
  );
  NAND _08070_ (
    .A(\memory[14][0] ),
    .B(_06002_),
    .Y(_06012_)
  );
  AND _08071_ (
    .A(_05403_),
    .B(_05454_),
    .Y(_06023_)
  );
  NAND _08072_ (
    .A(\memory[23][0] ),
    .B(_06023_),
    .Y(_06033_)
  );
  NOR _08073_ (
    .A(_05403_),
    .B(_05547_),
    .Y(_06043_)
  );
  NAND _08074_ (
    .A(\memory[2][0] ),
    .B(_06043_),
    .Y(_06054_)
  );
  AND _08075_ (
    .A(_05444_),
    .B(_05651_),
    .Y(_06064_)
  );
  NAND _08076_ (
    .A(\memory[15][0] ),
    .B(_06064_),
    .Y(_06074_)
  );
  AND _08077_ (
    .A(_05527_),
    .B(_05919_),
    .Y(_06085_)
  );
  NAND _08078_ (
    .A(\memory[16][0] ),
    .B(_06085_),
    .Y(_06095_)
  );
  AND _08079_ (
    .A(\op_addr[4] ),
    .B(_05382_),
    .Y(_06105_)
  );
  AND _08080_ (
    .A(\op_addr[0] ),
    .B(_06105_),
    .Y(_06116_)
  );
  NAND _08081_ (
    .A(\memory[1][0] ),
    .B(_06116_),
    .Y(_06126_)
  );
  NAND _08082_ (
    .A(_05506_),
    .B(_05775_),
    .Y(_06136_)
  );
  NOR _08083_ (
    .A(\op_addr[4] ),
    .B(_06136_),
    .Y(_06147_)
  );
  NAND _08084_ (
    .A(\memory[5][0] ),
    .B(_06147_),
    .Y(_06157_)
  );
  NOR _08085_ (
    .A(_05310_),
    .B(_06136_),
    .Y(_06167_)
  );
  NAND _08086_ (
    .A(\memory[21][0] ),
    .B(_06167_),
    .Y(_06178_)
  );
  AND _08087_ (
    .A(_05320_),
    .B(_06105_),
    .Y(_06188_)
  );
  NAND _08088_ (
    .A(\memory[0][0] ),
    .B(_06188_),
    .Y(_06198_)
  );
  AND _08089_ (
    .A(\op_addr[0] ),
    .B(_05392_),
    .Y(_06209_)
  );
  NAND _08090_ (
    .A(\memory[17][0] ),
    .B(_06209_),
    .Y(_06219_)
  );
  AND _08091_ (
    .A(_05775_),
    .B(_05868_),
    .Y(_06229_)
  );
  NAND _08092_ (
    .A(_05775_),
    .B(_05868_),
    .Y(_06240_)
  );
  AND _08093_ (
    .A(_05403_),
    .B(_06229_),
    .Y(_06250_)
  );
  NAND _08094_ (
    .A(\memory[25][0] ),
    .B(_06250_),
    .Y(_06260_)
  );
  AND _08095_ (
    .A(_05444_),
    .B(_05868_),
    .Y(_06271_)
  );
  NAND _08096_ (
    .A(_05444_),
    .B(_05868_),
    .Y(_06281_)
  );
  AND _08097_ (
    .A(_05403_),
    .B(_06271_),
    .Y(_06291_)
  );
  NAND _08098_ (
    .A(\memory[27][0] ),
    .B(_06291_),
    .Y(_06302_)
  );
  NOR _08099_ (
    .A(_05403_),
    .B(_06281_),
    .Y(_06312_)
  );
  NAND _08100_ (
    .A(\memory[11][0] ),
    .B(_06312_),
    .Y(_06322_)
  );
  AND _08101_ (
    .A(_05403_),
    .B(_05878_),
    .Y(_06333_)
  );
  NAND _08102_ (
    .A(\memory[26][0] ),
    .B(_06333_),
    .Y(_06343_)
  );
  NOR _08103_ (
    .A(_05403_),
    .B(_06240_),
    .Y(_06353_)
  );
  NAND _08104_ (
    .A(\memory[9][0] ),
    .B(_06353_),
    .Y(_06364_)
  );
  AND _08105_ (
    .A(_05868_),
    .B(_05950_),
    .Y(_06374_)
  );
  NAND _08106_ (
    .A(\memory[8][0] ),
    .B(_06374_),
    .Y(_06384_)
  );
  AND _08107_ (
    .A(_05868_),
    .B(_05919_),
    .Y(_06395_)
  );
  NAND _08108_ (
    .A(\memory[24][0] ),
    .B(_06395_),
    .Y(_06405_)
  );
  AND _08109_ (
    .A(_05795_),
    .B(_06074_),
    .Y(_06415_)
  );
  AND _08110_ (
    .A(_05816_),
    .B(_06415_),
    .Y(_06426_)
  );
  AND _08111_ (
    .A(_05857_),
    .B(_06426_),
    .Y(_06436_)
  );
  AND _08112_ (
    .A(_06033_),
    .B(_06054_),
    .Y(_06446_)
  );
  AND _08113_ (
    .A(_05837_),
    .B(_06012_),
    .Y(_06457_)
  );
  AND _08114_ (
    .A(_06446_),
    .B(_06457_),
    .Y(_06467_)
  );
  AND _08115_ (
    .A(_06436_),
    .B(_06467_),
    .Y(_06477_)
  );
  AND _08116_ (
    .A(_05568_),
    .B(_06157_),
    .Y(_06488_)
  );
  AND _08117_ (
    .A(_06126_),
    .B(_06198_),
    .Y(_06498_)
  );
  AND _08118_ (
    .A(_06178_),
    .B(_06219_),
    .Y(_06508_)
  );
  AND _08119_ (
    .A(_06498_),
    .B(_06508_),
    .Y(_06519_)
  );
  AND _08120_ (
    .A(_06488_),
    .B(_06519_),
    .Y(_06529_)
  );
  AND _08121_ (
    .A(_05940_),
    .B(_05971_),
    .Y(_06539_)
  );
  AND _08122_ (
    .A(_06529_),
    .B(_06539_),
    .Y(_06550_)
  );
  AND _08123_ (
    .A(_05609_),
    .B(_06405_),
    .Y(_06560_)
  );
  AND _08124_ (
    .A(_06302_),
    .B(_06364_),
    .Y(_06570_)
  );
  AND _08125_ (
    .A(_06560_),
    .B(_06570_),
    .Y(_06581_)
  );
  AND _08126_ (
    .A(_06550_),
    .B(_06581_),
    .Y(_06591_)
  );
  AND _08127_ (
    .A(_06477_),
    .B(_06591_),
    .Y(_06601_)
  );
  AND _08128_ (
    .A(_05671_),
    .B(_05744_),
    .Y(_06612_)
  );
  AND _08129_ (
    .A(_05702_),
    .B(_06612_),
    .Y(_06622_)
  );
  AND _08130_ (
    .A(_05485_),
    .B(_06622_),
    .Y(_06632_)
  );
  AND _08131_ (
    .A(_05909_),
    .B(_06384_),
    .Y(_06643_)
  );
  AND _08132_ (
    .A(_06260_),
    .B(_06343_),
    .Y(_06653_)
  );
  AND _08133_ (
    .A(_06643_),
    .B(_06653_),
    .Y(_06663_)
  );
  AND _08134_ (
    .A(_06095_),
    .B(_06322_),
    .Y(_06674_)
  );
  AND _08135_ (
    .A(_05764_),
    .B(_05992_),
    .Y(_06684_)
  );
  AND _08136_ (
    .A(_06674_),
    .B(_06684_),
    .Y(_06694_)
  );
  AND _08137_ (
    .A(_06663_),
    .B(_06694_),
    .Y(_06705_)
  );
  AND _08138_ (
    .A(_06632_),
    .B(_06705_),
    .Y(_06715_)
  );
  NAND _08139_ (
    .A(_06601_),
    .B(_06715_),
    .Y(\data_mem_o[16] )
  );
  NAND _08140_ (
    .A(\memory[22][1] ),
    .B(_05806_),
    .Y(_06735_)
  );
  NAND _08141_ (
    .A(\memory[3][1] ),
    .B(_05599_),
    .Y(_06745_)
  );
  NAND _08142_ (
    .A(\memory[12][1] ),
    .B(_05661_),
    .Y(_06755_)
  );
  NAND _08143_ (
    .A(\memory[29][1] ),
    .B(_05847_),
    .Y(_06766_)
  );
  NAND _08144_ (
    .A(\memory[23][1] ),
    .B(_06023_),
    .Y(_06776_)
  );
  NAND _08145_ (
    .A(\memory[13][1] ),
    .B(_05785_),
    .Y(_06786_)
  );
  NAND _08146_ (
    .A(\memory[19][1] ),
    .B(_05754_),
    .Y(_06797_)
  );
  NAND _08147_ (
    .A(\memory[31][1] ),
    .B(_05692_),
    .Y(_06807_)
  );
  NAND _08148_ (
    .A(\memory[2][1] ),
    .B(_06043_),
    .Y(_06817_)
  );
  NAND _08149_ (
    .A(\memory[6][1] ),
    .B(_05733_),
    .Y(_06828_)
  );
  NAND _08150_ (
    .A(\memory[30][1] ),
    .B(_05826_),
    .Y(_06838_)
  );
  NAND _08151_ (
    .A(\memory[11][1] ),
    .B(_06312_),
    .Y(_06848_)
  );
  NAND _08152_ (
    .A(\memory[27][1] ),
    .B(_06291_),
    .Y(_06859_)
  );
  NAND _08153_ (
    .A(\memory[25][1] ),
    .B(_06250_),
    .Y(_06869_)
  );
  NAND _08154_ (
    .A(\memory[24][1] ),
    .B(_06395_),
    .Y(_06879_)
  );
  NAND _08155_ (
    .A(\memory[14][1] ),
    .B(_06002_),
    .Y(_06890_)
  );
  NAND _08156_ (
    .A(\memory[15][1] ),
    .B(_06064_),
    .Y(_06900_)
  );
  AND _08157_ (
    .A(_06890_),
    .B(_06900_),
    .Y(_06910_)
  );
  NAND _08158_ (
    .A(\memory[7][1] ),
    .B(_05475_),
    .Y(_06921_)
  );
  NAND _08159_ (
    .A(\memory[18][1] ),
    .B(_05558_),
    .Y(_06931_)
  );
  NAND _08160_ (
    .A(\memory[9][1] ),
    .B(_06353_),
    .Y(_06941_)
  );
  NAND _08161_ (
    .A(\memory[0][1] ),
    .B(_06188_),
    .Y(_06952_)
  );
  NAND _08162_ (
    .A(\memory[17][1] ),
    .B(_06209_),
    .Y(_06962_)
  );
  NAND _08163_ (
    .A(\memory[1][1] ),
    .B(_06116_),
    .Y(_06972_)
  );
  NAND _08164_ (
    .A(\memory[5][1] ),
    .B(_06147_),
    .Y(_06983_)
  );
  NAND _08165_ (
    .A(\memory[21][1] ),
    .B(_06167_),
    .Y(_06993_)
  );
  NAND _08166_ (
    .A(\memory[8][1] ),
    .B(_06374_),
    .Y(_07003_)
  );
  NAND _08167_ (
    .A(\memory[20][1] ),
    .B(_05930_),
    .Y(_07014_)
  );
  NAND _08168_ (
    .A(\memory[10][1] ),
    .B(_05899_),
    .Y(_07024_)
  );
  NAND _08169_ (
    .A(\memory[26][1] ),
    .B(_06333_),
    .Y(_07034_)
  );
  NAND _08170_ (
    .A(\memory[4][1] ),
    .B(_05961_),
    .Y(_07045_)
  );
  NAND _08171_ (
    .A(\memory[16][1] ),
    .B(_06085_),
    .Y(_07055_)
  );
  NAND _08172_ (
    .A(\memory[28][1] ),
    .B(_05981_),
    .Y(_07065_)
  );
  AND _08173_ (
    .A(_06828_),
    .B(_06921_),
    .Y(_07076_)
  );
  AND _08174_ (
    .A(_06869_),
    .B(_07034_),
    .Y(_07086_)
  );
  AND _08175_ (
    .A(_06786_),
    .B(_06848_),
    .Y(_07096_)
  );
  AND _08176_ (
    .A(_07014_),
    .B(_07055_),
    .Y(_07107_)
  );
  AND _08177_ (
    .A(_07096_),
    .B(_07107_),
    .Y(_07117_)
  );
  AND _08178_ (
    .A(_06972_),
    .B(_07076_),
    .Y(_07127_)
  );
  AND _08179_ (
    .A(_06941_),
    .B(_07127_),
    .Y(_07138_)
  );
  AND _08180_ (
    .A(_07117_),
    .B(_07138_),
    .Y(_07148_)
  );
  AND _08181_ (
    .A(_06807_),
    .B(_06838_),
    .Y(_07158_)
  );
  AND _08182_ (
    .A(_06797_),
    .B(_07158_),
    .Y(_07169_)
  );
  AND _08183_ (
    .A(_07086_),
    .B(_07169_),
    .Y(_07179_)
  );
  AND _08184_ (
    .A(_06745_),
    .B(_06983_),
    .Y(_07189_)
  );
  AND _08185_ (
    .A(_06817_),
    .B(_07003_),
    .Y(_07200_)
  );
  AND _08186_ (
    .A(_07189_),
    .B(_07200_),
    .Y(_07210_)
  );
  AND _08187_ (
    .A(_07179_),
    .B(_07210_),
    .Y(_07220_)
  );
  AND _08188_ (
    .A(_07148_),
    .B(_07220_),
    .Y(_07231_)
  );
  AND _08189_ (
    .A(_06755_),
    .B(_07024_),
    .Y(_07241_)
  );
  AND _08190_ (
    .A(_06735_),
    .B(_06993_),
    .Y(_07251_)
  );
  AND _08191_ (
    .A(_07065_),
    .B(_07251_),
    .Y(_07262_)
  );
  AND _08192_ (
    .A(_07241_),
    .B(_07262_),
    .Y(_07272_)
  );
  AND _08193_ (
    .A(_06952_),
    .B(_07272_),
    .Y(_07282_)
  );
  AND _08194_ (
    .A(_06859_),
    .B(_06879_),
    .Y(_07293_)
  );
  AND _08195_ (
    .A(_06766_),
    .B(_07293_),
    .Y(_07303_)
  );
  AND _08196_ (
    .A(_06776_),
    .B(_06962_),
    .Y(_07313_)
  );
  AND _08197_ (
    .A(_06931_),
    .B(_07313_),
    .Y(_07324_)
  );
  AND _08198_ (
    .A(_06910_),
    .B(_07045_),
    .Y(_07334_)
  );
  AND _08199_ (
    .A(_07324_),
    .B(_07334_),
    .Y(_07345_)
  );
  AND _08200_ (
    .A(_07303_),
    .B(_07345_),
    .Y(_07356_)
  );
  AND _08201_ (
    .A(_07282_),
    .B(_07356_),
    .Y(_07367_)
  );
  NAND _08202_ (
    .A(_07231_),
    .B(_07367_),
    .Y(\data_mem_o[17] )
  );
  NAND _08203_ (
    .A(\memory[30][2] ),
    .B(_05826_),
    .Y(_07388_)
  );
  NAND _08204_ (
    .A(\memory[3][2] ),
    .B(_05599_),
    .Y(_07398_)
  );
  NAND _08205_ (
    .A(\memory[15][2] ),
    .B(_06064_),
    .Y(_07409_)
  );
  NAND _08206_ (
    .A(\memory[13][2] ),
    .B(_05785_),
    .Y(_07420_)
  );
  NAND _08207_ (
    .A(\memory[23][2] ),
    .B(_06023_),
    .Y(_07431_)
  );
  NAND _08208_ (
    .A(\memory[29][2] ),
    .B(_05847_),
    .Y(_07442_)
  );
  NAND _08209_ (
    .A(\memory[14][2] ),
    .B(_06002_),
    .Y(_07453_)
  );
  NAND _08210_ (
    .A(\memory[6][2] ),
    .B(_05733_),
    .Y(_07463_)
  );
  NAND _08211_ (
    .A(\memory[7][2] ),
    .B(_05475_),
    .Y(_07474_)
  );
  AND _08212_ (
    .A(_07463_),
    .B(_07474_),
    .Y(_07485_)
  );
  NAND _08213_ (
    .A(\memory[2][2] ),
    .B(_06043_),
    .Y(_07496_)
  );
  NAND _08214_ (
    .A(\memory[18][2] ),
    .B(_05558_),
    .Y(_07507_)
  );
  NAND _08215_ (
    .A(\memory[9][2] ),
    .B(_06353_),
    .Y(_07518_)
  );
  NAND _08216_ (
    .A(\memory[8][2] ),
    .B(_06374_),
    .Y(_07529_)
  );
  NAND _08217_ (
    .A(\memory[11][2] ),
    .B(_06312_),
    .Y(_07539_)
  );
  NAND _08218_ (
    .A(\memory[27][2] ),
    .B(_06291_),
    .Y(_07550_)
  );
  NAND _08219_ (
    .A(\memory[19][2] ),
    .B(_05754_),
    .Y(_07561_)
  );
  NAND _08220_ (
    .A(\memory[31][2] ),
    .B(_05692_),
    .Y(_07572_)
  );
  NAND _08221_ (
    .A(\memory[12][2] ),
    .B(_05661_),
    .Y(_07583_)
  );
  NAND _08222_ (
    .A(\memory[22][2] ),
    .B(_05806_),
    .Y(_07594_)
  );
  NAND _08223_ (
    .A(\memory[26][2] ),
    .B(_06333_),
    .Y(_07604_)
  );
  NAND _08224_ (
    .A(\memory[0][2] ),
    .B(_06188_),
    .Y(_07615_)
  );
  NAND _08225_ (
    .A(\memory[17][2] ),
    .B(_06209_),
    .Y(_07626_)
  );
  NAND _08226_ (
    .A(\memory[1][2] ),
    .B(_06116_),
    .Y(_07637_)
  );
  NAND _08227_ (
    .A(\memory[5][2] ),
    .B(_06147_),
    .Y(_07648_)
  );
  NAND _08228_ (
    .A(\memory[21][2] ),
    .B(_06167_),
    .Y(_07659_)
  );
  NAND _08229_ (
    .A(\memory[16][2] ),
    .B(_06085_),
    .Y(_07669_)
  );
  NAND _08230_ (
    .A(\memory[20][2] ),
    .B(_05930_),
    .Y(_07680_)
  );
  NAND _08231_ (
    .A(\memory[4][2] ),
    .B(_05961_),
    .Y(_07691_)
  );
  NAND _08232_ (
    .A(\memory[28][2] ),
    .B(_05981_),
    .Y(_07702_)
  );
  NAND _08233_ (
    .A(\memory[24][2] ),
    .B(_06395_),
    .Y(_07713_)
  );
  NAND _08234_ (
    .A(\memory[25][2] ),
    .B(_06250_),
    .Y(_07724_)
  );
  NAND _08235_ (
    .A(\memory[10][2] ),
    .B(_05899_),
    .Y(_07734_)
  );
  AND _08236_ (
    .A(_07604_),
    .B(_07724_),
    .Y(_07745_)
  );
  AND _08237_ (
    .A(_07420_),
    .B(_07539_),
    .Y(_07756_)
  );
  AND _08238_ (
    .A(_07669_),
    .B(_07680_),
    .Y(_07767_)
  );
  AND _08239_ (
    .A(_07756_),
    .B(_07767_),
    .Y(_07778_)
  );
  AND _08240_ (
    .A(_07485_),
    .B(_07637_),
    .Y(_07789_)
  );
  AND _08241_ (
    .A(_07518_),
    .B(_07789_),
    .Y(_07800_)
  );
  AND _08242_ (
    .A(_07778_),
    .B(_07800_),
    .Y(_07810_)
  );
  AND _08243_ (
    .A(_07388_),
    .B(_07572_),
    .Y(_07821_)
  );
  AND _08244_ (
    .A(_07561_),
    .B(_07821_),
    .Y(_07832_)
  );
  AND _08245_ (
    .A(_07745_),
    .B(_07832_),
    .Y(_07843_)
  );
  AND _08246_ (
    .A(_07398_),
    .B(_07648_),
    .Y(_07854_)
  );
  AND _08247_ (
    .A(_07496_),
    .B(_07529_),
    .Y(_07865_)
  );
  AND _08248_ (
    .A(_07854_),
    .B(_07865_),
    .Y(_07871_)
  );
  AND _08249_ (
    .A(_07843_),
    .B(_07871_),
    .Y(_07872_)
  );
  AND _08250_ (
    .A(_07810_),
    .B(_07872_),
    .Y(_07873_)
  );
  AND _08251_ (
    .A(_07583_),
    .B(_07734_),
    .Y(_07874_)
  );
  AND _08252_ (
    .A(_07594_),
    .B(_07659_),
    .Y(_07875_)
  );
  AND _08253_ (
    .A(_07702_),
    .B(_07875_),
    .Y(_07876_)
  );
  AND _08254_ (
    .A(_07874_),
    .B(_07876_),
    .Y(_07877_)
  );
  AND _08255_ (
    .A(_07615_),
    .B(_07877_),
    .Y(_07878_)
  );
  AND _08256_ (
    .A(_07550_),
    .B(_07713_),
    .Y(_07879_)
  );
  AND _08257_ (
    .A(_07442_),
    .B(_07879_),
    .Y(_07880_)
  );
  AND _08258_ (
    .A(_07431_),
    .B(_07626_),
    .Y(_07881_)
  );
  AND _08259_ (
    .A(_07507_),
    .B(_07881_),
    .Y(_07882_)
  );
  AND _08260_ (
    .A(_07409_),
    .B(_07453_),
    .Y(_07883_)
  );
  AND _08261_ (
    .A(_07691_),
    .B(_07883_),
    .Y(_07884_)
  );
  AND _08262_ (
    .A(_07882_),
    .B(_07884_),
    .Y(_07885_)
  );
  AND _08263_ (
    .A(_07880_),
    .B(_07885_),
    .Y(_07886_)
  );
  AND _08264_ (
    .A(_07878_),
    .B(_07886_),
    .Y(_07887_)
  );
  NAND _08265_ (
    .A(_07873_),
    .B(_07887_),
    .Y(\data_mem_o[18] )
  );
  NAND _08266_ (
    .A(\memory[6][3] ),
    .B(_05733_),
    .Y(_07888_)
  );
  NAND _08267_ (
    .A(\memory[19][3] ),
    .B(_05754_),
    .Y(_07889_)
  );
  NAND _08268_ (
    .A(\memory[3][3] ),
    .B(_05599_),
    .Y(_07890_)
  );
  NAND _08269_ (
    .A(\memory[30][3] ),
    .B(_05826_),
    .Y(_07891_)
  );
  NAND _08270_ (
    .A(\memory[22][3] ),
    .B(_05806_),
    .Y(_07892_)
  );
  NAND _08271_ (
    .A(\memory[23][3] ),
    .B(_06023_),
    .Y(_07893_)
  );
  NAND _08272_ (
    .A(\memory[18][3] ),
    .B(_05558_),
    .Y(_07894_)
  );
  NAND _08273_ (
    .A(\memory[12][3] ),
    .B(_05661_),
    .Y(_07895_)
  );
  NAND _08274_ (
    .A(\memory[31][3] ),
    .B(_05692_),
    .Y(_07896_)
  );
  NAND _08275_ (
    .A(\memory[7][3] ),
    .B(_05475_),
    .Y(_07897_)
  );
  NAND _08276_ (
    .A(\memory[29][3] ),
    .B(_05847_),
    .Y(_07898_)
  );
  NAND _08277_ (
    .A(\memory[10][3] ),
    .B(_05899_),
    .Y(_07899_)
  );
  NAND _08278_ (
    .A(\memory[9][3] ),
    .B(_06353_),
    .Y(_07900_)
  );
  NAND _08279_ (
    .A(\memory[28][3] ),
    .B(_05981_),
    .Y(_07901_)
  );
  NAND _08280_ (
    .A(\memory[24][3] ),
    .B(_06395_),
    .Y(_07902_)
  );
  NAND _08281_ (
    .A(\memory[15][3] ),
    .B(_06064_),
    .Y(_07903_)
  );
  NAND _08282_ (
    .A(\memory[14][3] ),
    .B(_06002_),
    .Y(_07904_)
  );
  AND _08283_ (
    .A(_07903_),
    .B(_07904_),
    .Y(_07905_)
  );
  NAND _08284_ (
    .A(\memory[13][3] ),
    .B(_05785_),
    .Y(_07906_)
  );
  NAND _08285_ (
    .A(\memory[2][3] ),
    .B(_06043_),
    .Y(_07907_)
  );
  NAND _08286_ (
    .A(\memory[26][3] ),
    .B(_06333_),
    .Y(_07908_)
  );
  NAND _08287_ (
    .A(\memory[17][3] ),
    .B(_06209_),
    .Y(_07909_)
  );
  NAND _08288_ (
    .A(\memory[0][3] ),
    .B(_06188_),
    .Y(_07910_)
  );
  NAND _08289_ (
    .A(\memory[1][3] ),
    .B(_06116_),
    .Y(_07911_)
  );
  NAND _08290_ (
    .A(\memory[21][3] ),
    .B(_06167_),
    .Y(_07912_)
  );
  NAND _08291_ (
    .A(\memory[5][3] ),
    .B(_06147_),
    .Y(_07913_)
  );
  NAND _08292_ (
    .A(\memory[11][3] ),
    .B(_06312_),
    .Y(_07914_)
  );
  NAND _08293_ (
    .A(\memory[27][3] ),
    .B(_06291_),
    .Y(_07915_)
  );
  NAND _08294_ (
    .A(\memory[8][3] ),
    .B(_06374_),
    .Y(_07916_)
  );
  NAND _08295_ (
    .A(\memory[25][3] ),
    .B(_06250_),
    .Y(_07917_)
  );
  NAND _08296_ (
    .A(\memory[16][3] ),
    .B(_06085_),
    .Y(_07918_)
  );
  NAND _08297_ (
    .A(\memory[20][3] ),
    .B(_05930_),
    .Y(_07919_)
  );
  NAND _08298_ (
    .A(\memory[4][3] ),
    .B(_05961_),
    .Y(_07920_)
  );
  AND _08299_ (
    .A(_07914_),
    .B(_07918_),
    .Y(_07921_)
  );
  AND _08300_ (
    .A(_07888_),
    .B(_07897_),
    .Y(_07922_)
  );
  AND _08301_ (
    .A(_07893_),
    .B(_07912_),
    .Y(_07923_)
  );
  AND _08302_ (
    .A(_07911_),
    .B(_07923_),
    .Y(_07924_)
  );
  AND _08303_ (
    .A(_07922_),
    .B(_07924_),
    .Y(_07925_)
  );
  AND _08304_ (
    .A(_07895_),
    .B(_07899_),
    .Y(_07926_)
  );
  AND _08305_ (
    .A(_07915_),
    .B(_07926_),
    .Y(_07927_)
  );
  AND _08306_ (
    .A(_07925_),
    .B(_07927_),
    .Y(_07928_)
  );
  AND _08307_ (
    .A(_07906_),
    .B(_07919_),
    .Y(_07929_)
  );
  AND _08308_ (
    .A(_07928_),
    .B(_07929_),
    .Y(_07930_)
  );
  AND _08309_ (
    .A(_07901_),
    .B(_07917_),
    .Y(_07931_)
  );
  AND _08310_ (
    .A(_07891_),
    .B(_07898_),
    .Y(_07932_)
  );
  AND _08311_ (
    .A(_07900_),
    .B(_07932_),
    .Y(_07933_)
  );
  AND _08312_ (
    .A(_07896_),
    .B(_07933_),
    .Y(_07934_)
  );
  AND _08313_ (
    .A(_07894_),
    .B(_07902_),
    .Y(_07935_)
  );
  AND _08314_ (
    .A(_07889_),
    .B(_07935_),
    .Y(_07936_)
  );
  AND _08315_ (
    .A(_07934_),
    .B(_07936_),
    .Y(_07937_)
  );
  AND _08316_ (
    .A(_07931_),
    .B(_07937_),
    .Y(_07938_)
  );
  AND _08317_ (
    .A(_07930_),
    .B(_07938_),
    .Y(_07939_)
  );
  AND _08318_ (
    .A(_07890_),
    .B(_07907_),
    .Y(_07940_)
  );
  AND _08319_ (
    .A(_07921_),
    .B(_07940_),
    .Y(_07941_)
  );
  AND _08320_ (
    .A(_07892_),
    .B(_07909_),
    .Y(_07942_)
  );
  AND _08321_ (
    .A(_07913_),
    .B(_07916_),
    .Y(_07943_)
  );
  AND _08322_ (
    .A(_07942_),
    .B(_07943_),
    .Y(_07944_)
  );
  AND _08323_ (
    .A(_07908_),
    .B(_07910_),
    .Y(_07945_)
  );
  AND _08324_ (
    .A(_07905_),
    .B(_07920_),
    .Y(_07946_)
  );
  AND _08325_ (
    .A(_07945_),
    .B(_07946_),
    .Y(_07947_)
  );
  AND _08326_ (
    .A(_07944_),
    .B(_07947_),
    .Y(_07948_)
  );
  AND _08327_ (
    .A(_07941_),
    .B(_07948_),
    .Y(_07949_)
  );
  NAND _08328_ (
    .A(_07939_),
    .B(_07949_),
    .Y(\data_mem_o[19] )
  );
  NAND _08329_ (
    .A(\memory[2][4] ),
    .B(_06043_),
    .Y(_07950_)
  );
  NAND _08330_ (
    .A(\memory[7][4] ),
    .B(_05475_),
    .Y(_07951_)
  );
  NAND _08331_ (
    .A(\memory[29][4] ),
    .B(_05847_),
    .Y(_07952_)
  );
  AND _08332_ (
    .A(_07951_),
    .B(_07952_),
    .Y(_07953_)
  );
  AND _08333_ (
    .A(_07950_),
    .B(_07953_),
    .Y(_07954_)
  );
  NAND _08334_ (
    .A(\memory[19][4] ),
    .B(_05754_),
    .Y(_07955_)
  );
  NAND _08335_ (
    .A(\memory[3][4] ),
    .B(_05599_),
    .Y(_07956_)
  );
  AND _08336_ (
    .A(_07955_),
    .B(_07956_),
    .Y(_07957_)
  );
  NAND _08337_ (
    .A(\memory[12][4] ),
    .B(_05661_),
    .Y(_07958_)
  );
  NAND _08338_ (
    .A(\memory[13][4] ),
    .B(_05785_),
    .Y(_07959_)
  );
  AND _08339_ (
    .A(_07958_),
    .B(_07959_),
    .Y(_07960_)
  );
  AND _08340_ (
    .A(_07957_),
    .B(_07960_),
    .Y(_07961_)
  );
  NAND _08341_ (
    .A(\memory[31][4] ),
    .B(_05692_),
    .Y(_07962_)
  );
  NAND _08342_ (
    .A(\memory[30][4] ),
    .B(_05826_),
    .Y(_07963_)
  );
  AND _08343_ (
    .A(_07962_),
    .B(_07963_),
    .Y(_07964_)
  );
  NAND _08344_ (
    .A(\memory[14][4] ),
    .B(_06002_),
    .Y(_07965_)
  );
  NAND _08345_ (
    .A(\memory[15][4] ),
    .B(_06064_),
    .Y(_07966_)
  );
  AND _08346_ (
    .A(_07965_),
    .B(_07966_),
    .Y(_07967_)
  );
  AND _08347_ (
    .A(_07964_),
    .B(_07967_),
    .Y(_07968_)
  );
  AND _08348_ (
    .A(_07961_),
    .B(_07968_),
    .Y(_07969_)
  );
  AND _08349_ (
    .A(_07954_),
    .B(_07969_),
    .Y(_07970_)
  );
  NAND _08350_ (
    .A(\memory[9][4] ),
    .B(_06353_),
    .Y(_07971_)
  );
  NAND _08351_ (
    .A(\memory[27][4] ),
    .B(_06291_),
    .Y(_07972_)
  );
  AND _08352_ (
    .A(_07971_),
    .B(_07972_),
    .Y(_07973_)
  );
  NAND _08353_ (
    .A(\memory[16][4] ),
    .B(_06085_),
    .Y(_07974_)
  );
  NAND _08354_ (
    .A(\memory[8][4] ),
    .B(_06374_),
    .Y(_07975_)
  );
  AND _08355_ (
    .A(_07974_),
    .B(_07975_),
    .Y(_07976_)
  );
  AND _08356_ (
    .A(_07973_),
    .B(_07976_),
    .Y(_07977_)
  );
  NAND _08357_ (
    .A(\memory[18][4] ),
    .B(_05558_),
    .Y(_07978_)
  );
  NAND _08358_ (
    .A(\memory[23][4] ),
    .B(_06023_),
    .Y(_07979_)
  );
  AND _08359_ (
    .A(_07978_),
    .B(_07979_),
    .Y(_07980_)
  );
  NAND _08360_ (
    .A(\memory[22][4] ),
    .B(_05806_),
    .Y(_07981_)
  );
  NAND _08361_ (
    .A(\memory[6][4] ),
    .B(_05733_),
    .Y(_07982_)
  );
  AND _08362_ (
    .A(_07981_),
    .B(_07982_),
    .Y(_07983_)
  );
  AND _08363_ (
    .A(_07980_),
    .B(_07983_),
    .Y(_07984_)
  );
  NAND _08364_ (
    .A(\memory[24][4] ),
    .B(_06395_),
    .Y(_07985_)
  );
  NAND _08365_ (
    .A(\memory[17][4] ),
    .B(_06209_),
    .Y(_07986_)
  );
  NAND _08366_ (
    .A(\memory[21][4] ),
    .B(_06167_),
    .Y(_07987_)
  );
  NAND _08367_ (
    .A(\memory[5][4] ),
    .B(_06147_),
    .Y(_07988_)
  );
  AND _08368_ (
    .A(_07987_),
    .B(_07988_),
    .Y(_07989_)
  );
  AND _08369_ (
    .A(_07986_),
    .B(_07989_),
    .Y(_07990_)
  );
  NAND _08370_ (
    .A(\memory[0][4] ),
    .B(_06188_),
    .Y(_07991_)
  );
  NAND _08371_ (
    .A(\memory[1][4] ),
    .B(_06116_),
    .Y(_07992_)
  );
  AND _08372_ (
    .A(_07991_),
    .B(_07992_),
    .Y(_07993_)
  );
  AND _08373_ (
    .A(_07990_),
    .B(_07993_),
    .Y(_07994_)
  );
  AND _08374_ (
    .A(_07985_),
    .B(_07994_),
    .Y(_07995_)
  );
  AND _08375_ (
    .A(_07984_),
    .B(_07995_),
    .Y(_07996_)
  );
  AND _08376_ (
    .A(_07977_),
    .B(_07996_),
    .Y(_07997_)
  );
  NAND _08377_ (
    .A(\memory[20][4] ),
    .B(_05930_),
    .Y(_07998_)
  );
  NAND _08378_ (
    .A(\memory[28][4] ),
    .B(_05981_),
    .Y(_07999_)
  );
  NAND _08379_ (
    .A(\memory[11][4] ),
    .B(_06312_),
    .Y(_08000_)
  );
  AND _08380_ (
    .A(_07999_),
    .B(_08000_),
    .Y(_00256_)
  );
  AND _08381_ (
    .A(_07998_),
    .B(_00256_),
    .Y(_00257_)
  );
  NAND _08382_ (
    .A(\memory[25][4] ),
    .B(_06250_),
    .Y(_00258_)
  );
  NAND _08383_ (
    .A(\memory[26][4] ),
    .B(_06333_),
    .Y(_00259_)
  );
  AND _08384_ (
    .A(_00258_),
    .B(_00259_),
    .Y(_00260_)
  );
  NAND _08385_ (
    .A(\memory[10][4] ),
    .B(_05899_),
    .Y(_00261_)
  );
  NAND _08386_ (
    .A(\memory[4][4] ),
    .B(_05961_),
    .Y(_00262_)
  );
  AND _08387_ (
    .A(_00261_),
    .B(_00262_),
    .Y(_00263_)
  );
  AND _08388_ (
    .A(_00260_),
    .B(_00263_),
    .Y(_00264_)
  );
  AND _08389_ (
    .A(_00257_),
    .B(_00264_),
    .Y(_00265_)
  );
  AND _08390_ (
    .A(_07997_),
    .B(_00265_),
    .Y(_00266_)
  );
  NAND _08391_ (
    .A(_07970_),
    .B(_00266_),
    .Y(\data_mem_o[20] )
  );
  NAND _08392_ (
    .A(\memory[22][5] ),
    .B(_05806_),
    .Y(_00267_)
  );
  NAND _08393_ (
    .A(\memory[3][5] ),
    .B(_05599_),
    .Y(_00268_)
  );
  NAND _08394_ (
    .A(\memory[12][5] ),
    .B(_05661_),
    .Y(_00269_)
  );
  NAND _08395_ (
    .A(\memory[29][5] ),
    .B(_05847_),
    .Y(_00270_)
  );
  NAND _08396_ (
    .A(\memory[23][5] ),
    .B(_06023_),
    .Y(_00271_)
  );
  NAND _08397_ (
    .A(\memory[13][5] ),
    .B(_05785_),
    .Y(_00272_)
  );
  NAND _08398_ (
    .A(\memory[19][5] ),
    .B(_05754_),
    .Y(_00273_)
  );
  NAND _08399_ (
    .A(\memory[31][5] ),
    .B(_05692_),
    .Y(_00274_)
  );
  NAND _08400_ (
    .A(\memory[2][5] ),
    .B(_06043_),
    .Y(_00275_)
  );
  NAND _08401_ (
    .A(\memory[6][5] ),
    .B(_05733_),
    .Y(_00276_)
  );
  NAND _08402_ (
    .A(\memory[30][5] ),
    .B(_05826_),
    .Y(_00277_)
  );
  NAND _08403_ (
    .A(\memory[11][5] ),
    .B(_06312_),
    .Y(_00278_)
  );
  NAND _08404_ (
    .A(\memory[27][5] ),
    .B(_06291_),
    .Y(_00279_)
  );
  NAND _08405_ (
    .A(\memory[25][5] ),
    .B(_06250_),
    .Y(_00280_)
  );
  NAND _08406_ (
    .A(\memory[24][5] ),
    .B(_06395_),
    .Y(_00281_)
  );
  NAND _08407_ (
    .A(\memory[14][5] ),
    .B(_06002_),
    .Y(_00282_)
  );
  NAND _08408_ (
    .A(\memory[15][5] ),
    .B(_06064_),
    .Y(_00283_)
  );
  AND _08409_ (
    .A(_00282_),
    .B(_00283_),
    .Y(_00284_)
  );
  NAND _08410_ (
    .A(\memory[7][5] ),
    .B(_05475_),
    .Y(_00285_)
  );
  NAND _08411_ (
    .A(\memory[18][5] ),
    .B(_05558_),
    .Y(_00286_)
  );
  NAND _08412_ (
    .A(\memory[9][5] ),
    .B(_06353_),
    .Y(_00287_)
  );
  NAND _08413_ (
    .A(\memory[0][5] ),
    .B(_06188_),
    .Y(_00288_)
  );
  NAND _08414_ (
    .A(\memory[17][5] ),
    .B(_06209_),
    .Y(_00289_)
  );
  NAND _08415_ (
    .A(\memory[1][5] ),
    .B(_06116_),
    .Y(_00290_)
  );
  NAND _08416_ (
    .A(\memory[5][5] ),
    .B(_06147_),
    .Y(_00291_)
  );
  NAND _08417_ (
    .A(\memory[21][5] ),
    .B(_06167_),
    .Y(_00292_)
  );
  NAND _08418_ (
    .A(\memory[8][5] ),
    .B(_06374_),
    .Y(_00293_)
  );
  NAND _08419_ (
    .A(\memory[20][5] ),
    .B(_05930_),
    .Y(_00294_)
  );
  NAND _08420_ (
    .A(\memory[10][5] ),
    .B(_05899_),
    .Y(_00295_)
  );
  NAND _08421_ (
    .A(\memory[26][5] ),
    .B(_06333_),
    .Y(_00296_)
  );
  NAND _08422_ (
    .A(\memory[4][5] ),
    .B(_05961_),
    .Y(_00297_)
  );
  NAND _08423_ (
    .A(\memory[16][5] ),
    .B(_06085_),
    .Y(_00298_)
  );
  NAND _08424_ (
    .A(\memory[28][5] ),
    .B(_05981_),
    .Y(_00299_)
  );
  AND _08425_ (
    .A(_00276_),
    .B(_00285_),
    .Y(_00300_)
  );
  AND _08426_ (
    .A(_00280_),
    .B(_00296_),
    .Y(_00301_)
  );
  AND _08427_ (
    .A(_00272_),
    .B(_00278_),
    .Y(_00302_)
  );
  AND _08428_ (
    .A(_00294_),
    .B(_00298_),
    .Y(_00303_)
  );
  AND _08429_ (
    .A(_00302_),
    .B(_00303_),
    .Y(_00304_)
  );
  AND _08430_ (
    .A(_00290_),
    .B(_00300_),
    .Y(_00305_)
  );
  AND _08431_ (
    .A(_00287_),
    .B(_00305_),
    .Y(_00306_)
  );
  AND _08432_ (
    .A(_00304_),
    .B(_00306_),
    .Y(_00307_)
  );
  AND _08433_ (
    .A(_00274_),
    .B(_00277_),
    .Y(_00308_)
  );
  AND _08434_ (
    .A(_00273_),
    .B(_00308_),
    .Y(_00309_)
  );
  AND _08435_ (
    .A(_00301_),
    .B(_00309_),
    .Y(_00310_)
  );
  AND _08436_ (
    .A(_00268_),
    .B(_00291_),
    .Y(_00311_)
  );
  AND _08437_ (
    .A(_00275_),
    .B(_00293_),
    .Y(_00312_)
  );
  AND _08438_ (
    .A(_00311_),
    .B(_00312_),
    .Y(_00313_)
  );
  AND _08439_ (
    .A(_00310_),
    .B(_00313_),
    .Y(_00314_)
  );
  AND _08440_ (
    .A(_00307_),
    .B(_00314_),
    .Y(_00315_)
  );
  AND _08441_ (
    .A(_00269_),
    .B(_00295_),
    .Y(_00316_)
  );
  AND _08442_ (
    .A(_00267_),
    .B(_00292_),
    .Y(_00317_)
  );
  AND _08443_ (
    .A(_00299_),
    .B(_00317_),
    .Y(_00318_)
  );
  AND _08444_ (
    .A(_00316_),
    .B(_00318_),
    .Y(_00319_)
  );
  AND _08445_ (
    .A(_00288_),
    .B(_00319_),
    .Y(_00320_)
  );
  AND _08446_ (
    .A(_00279_),
    .B(_00281_),
    .Y(_00321_)
  );
  AND _08447_ (
    .A(_00270_),
    .B(_00321_),
    .Y(_00322_)
  );
  AND _08448_ (
    .A(_00271_),
    .B(_00289_),
    .Y(_00323_)
  );
  AND _08449_ (
    .A(_00286_),
    .B(_00323_),
    .Y(_00324_)
  );
  AND _08450_ (
    .A(_00284_),
    .B(_00297_),
    .Y(_00325_)
  );
  AND _08451_ (
    .A(_00324_),
    .B(_00325_),
    .Y(_00326_)
  );
  AND _08452_ (
    .A(_00322_),
    .B(_00326_),
    .Y(_00327_)
  );
  AND _08453_ (
    .A(_00320_),
    .B(_00327_),
    .Y(_00328_)
  );
  NAND _08454_ (
    .A(_00315_),
    .B(_00328_),
    .Y(\data_mem_o[21] )
  );
  NAND _08455_ (
    .A(\memory[7][6] ),
    .B(_05475_),
    .Y(_00329_)
  );
  NAND _08456_ (
    .A(\memory[14][6] ),
    .B(_06002_),
    .Y(_00330_)
  );
  NAND _08457_ (
    .A(\memory[15][6] ),
    .B(_06064_),
    .Y(_00331_)
  );
  NAND _08458_ (
    .A(\memory[29][6] ),
    .B(_05847_),
    .Y(_00332_)
  );
  NAND _08459_ (
    .A(\memory[19][6] ),
    .B(_05754_),
    .Y(_00333_)
  );
  NAND _08460_ (
    .A(\memory[3][6] ),
    .B(_05599_),
    .Y(_00334_)
  );
  NAND _08461_ (
    .A(\memory[2][6] ),
    .B(_06043_),
    .Y(_00335_)
  );
  NAND _08462_ (
    .A(\memory[13][6] ),
    .B(_05785_),
    .Y(_00336_)
  );
  NAND _08463_ (
    .A(\memory[18][6] ),
    .B(_05558_),
    .Y(_00337_)
  );
  NAND _08464_ (
    .A(\memory[30][6] ),
    .B(_05826_),
    .Y(_00338_)
  );
  NAND _08465_ (
    .A(\memory[31][6] ),
    .B(_05692_),
    .Y(_00339_)
  );
  NAND _08466_ (
    .A(\memory[4][6] ),
    .B(_05961_),
    .Y(_00340_)
  );
  NAND _08467_ (
    .A(\memory[8][6] ),
    .B(_06374_),
    .Y(_00341_)
  );
  NAND _08468_ (
    .A(\memory[9][6] ),
    .B(_06353_),
    .Y(_00342_)
  );
  NAND _08469_ (
    .A(\memory[25][6] ),
    .B(_06250_),
    .Y(_00343_)
  );
  NAND _08470_ (
    .A(\memory[12][6] ),
    .B(_05661_),
    .Y(_00344_)
  );
  NAND _08471_ (
    .A(\memory[6][6] ),
    .B(_05733_),
    .Y(_00345_)
  );
  NAND _08472_ (
    .A(\memory[22][6] ),
    .B(_05806_),
    .Y(_00346_)
  );
  NAND _08473_ (
    .A(\memory[23][6] ),
    .B(_06023_),
    .Y(_00347_)
  );
  NAND _08474_ (
    .A(\memory[16][6] ),
    .B(_06085_),
    .Y(_00348_)
  );
  NAND _08475_ (
    .A(\memory[17][6] ),
    .B(_06209_),
    .Y(_00349_)
  );
  NAND _08476_ (
    .A(\memory[21][6] ),
    .B(_06167_),
    .Y(_00350_)
  );
  NAND _08477_ (
    .A(\memory[5][6] ),
    .B(_06147_),
    .Y(_00351_)
  );
  NAND _08478_ (
    .A(\memory[1][6] ),
    .B(_06116_),
    .Y(_00352_)
  );
  NAND _08479_ (
    .A(\memory[0][6] ),
    .B(_06188_),
    .Y(_00353_)
  );
  NAND _08480_ (
    .A(\memory[27][6] ),
    .B(_06291_),
    .Y(_00354_)
  );
  NAND _08481_ (
    .A(\memory[10][6] ),
    .B(_05899_),
    .Y(_00355_)
  );
  NAND _08482_ (
    .A(\memory[26][6] ),
    .B(_06333_),
    .Y(_00356_)
  );
  NAND _08483_ (
    .A(\memory[20][6] ),
    .B(_05930_),
    .Y(_00357_)
  );
  NAND _08484_ (
    .A(\memory[28][6] ),
    .B(_05981_),
    .Y(_00358_)
  );
  NAND _08485_ (
    .A(\memory[24][6] ),
    .B(_06395_),
    .Y(_00359_)
  );
  NAND _08486_ (
    .A(\memory[11][6] ),
    .B(_06312_),
    .Y(_00360_)
  );
  AND _08487_ (
    .A(_00337_),
    .B(_00347_),
    .Y(_00361_)
  );
  AND _08488_ (
    .A(_00330_),
    .B(_00334_),
    .Y(_00362_)
  );
  AND _08489_ (
    .A(_00344_),
    .B(_00355_),
    .Y(_00363_)
  );
  AND _08490_ (
    .A(_00345_),
    .B(_00352_),
    .Y(_00364_)
  );
  AND _08491_ (
    .A(_00363_),
    .B(_00364_),
    .Y(_00365_)
  );
  AND _08492_ (
    .A(_00362_),
    .B(_00365_),
    .Y(_00366_)
  );
  AND _08493_ (
    .A(_00346_),
    .B(_00349_),
    .Y(_00367_)
  );
  AND _08494_ (
    .A(_00342_),
    .B(_00367_),
    .Y(_00368_)
  );
  AND _08495_ (
    .A(_00350_),
    .B(_00368_),
    .Y(_00369_)
  );
  AND _08496_ (
    .A(_00357_),
    .B(_00369_),
    .Y(_00370_)
  );
  AND _08497_ (
    .A(_00366_),
    .B(_00370_),
    .Y(_00371_)
  );
  AND _08498_ (
    .A(_00335_),
    .B(_00340_),
    .Y(_00372_)
  );
  AND _08499_ (
    .A(_00331_),
    .B(_00372_),
    .Y(_00373_)
  );
  AND _08500_ (
    .A(_00341_),
    .B(_00351_),
    .Y(_00374_)
  );
  AND _08501_ (
    .A(_00329_),
    .B(_00374_),
    .Y(_00375_)
  );
  AND _08502_ (
    .A(_00373_),
    .B(_00375_),
    .Y(_00376_)
  );
  AND _08503_ (
    .A(_00338_),
    .B(_00343_),
    .Y(_00377_)
  );
  AND _08504_ (
    .A(_00354_),
    .B(_00356_),
    .Y(_00378_)
  );
  AND _08505_ (
    .A(_00332_),
    .B(_00378_),
    .Y(_00379_)
  );
  AND _08506_ (
    .A(_00377_),
    .B(_00379_),
    .Y(_00380_)
  );
  AND _08507_ (
    .A(_00376_),
    .B(_00380_),
    .Y(_00381_)
  );
  AND _08508_ (
    .A(_00371_),
    .B(_00381_),
    .Y(_00382_)
  );
  AND _08509_ (
    .A(_00339_),
    .B(_00358_),
    .Y(_00383_)
  );
  AND _08510_ (
    .A(_00333_),
    .B(_00348_),
    .Y(_00384_)
  );
  AND _08511_ (
    .A(_00383_),
    .B(_00384_),
    .Y(_00385_)
  );
  AND _08512_ (
    .A(_00336_),
    .B(_00360_),
    .Y(_00386_)
  );
  AND _08513_ (
    .A(_00353_),
    .B(_00361_),
    .Y(_00387_)
  );
  AND _08514_ (
    .A(_00386_),
    .B(_00387_),
    .Y(_00388_)
  );
  AND _08515_ (
    .A(_00385_),
    .B(_00388_),
    .Y(_00389_)
  );
  AND _08516_ (
    .A(_00359_),
    .B(_00389_),
    .Y(_00390_)
  );
  NAND _08517_ (
    .A(_00382_),
    .B(_00390_),
    .Y(\data_mem_o[22] )
  );
  NAND _08518_ (
    .A(\memory[22][7] ),
    .B(_05806_),
    .Y(_00391_)
  );
  NAND _08519_ (
    .A(\memory[3][7] ),
    .B(_05599_),
    .Y(_00392_)
  );
  NAND _08520_ (
    .A(\memory[12][7] ),
    .B(_05661_),
    .Y(_00393_)
  );
  NAND _08521_ (
    .A(\memory[29][7] ),
    .B(_05847_),
    .Y(_00394_)
  );
  NAND _08522_ (
    .A(\memory[23][7] ),
    .B(_06023_),
    .Y(_00395_)
  );
  NAND _08523_ (
    .A(\memory[13][7] ),
    .B(_05785_),
    .Y(_00396_)
  );
  NAND _08524_ (
    .A(\memory[19][7] ),
    .B(_05754_),
    .Y(_00397_)
  );
  NAND _08525_ (
    .A(\memory[31][7] ),
    .B(_05692_),
    .Y(_00398_)
  );
  NAND _08526_ (
    .A(\memory[2][7] ),
    .B(_06043_),
    .Y(_00399_)
  );
  NAND _08527_ (
    .A(\memory[6][7] ),
    .B(_05733_),
    .Y(_00400_)
  );
  NAND _08528_ (
    .A(\memory[30][7] ),
    .B(_05826_),
    .Y(_00401_)
  );
  NAND _08529_ (
    .A(\memory[11][7] ),
    .B(_06312_),
    .Y(_00402_)
  );
  NAND _08530_ (
    .A(\memory[27][7] ),
    .B(_06291_),
    .Y(_00403_)
  );
  NAND _08531_ (
    .A(\memory[25][7] ),
    .B(_06250_),
    .Y(_00404_)
  );
  NAND _08532_ (
    .A(\memory[24][7] ),
    .B(_06395_),
    .Y(_00405_)
  );
  NAND _08533_ (
    .A(\memory[14][7] ),
    .B(_06002_),
    .Y(_00406_)
  );
  NAND _08534_ (
    .A(\memory[15][7] ),
    .B(_06064_),
    .Y(_00407_)
  );
  AND _08535_ (
    .A(_00406_),
    .B(_00407_),
    .Y(_00408_)
  );
  NAND _08536_ (
    .A(\memory[7][7] ),
    .B(_05475_),
    .Y(_00409_)
  );
  NAND _08537_ (
    .A(\memory[18][7] ),
    .B(_05558_),
    .Y(_00410_)
  );
  NAND _08538_ (
    .A(\memory[9][7] ),
    .B(_06353_),
    .Y(_00411_)
  );
  NAND _08539_ (
    .A(\memory[0][7] ),
    .B(_06188_),
    .Y(_00412_)
  );
  NAND _08540_ (
    .A(\memory[17][7] ),
    .B(_06209_),
    .Y(_00413_)
  );
  NAND _08541_ (
    .A(\memory[1][7] ),
    .B(_06116_),
    .Y(_00414_)
  );
  NAND _08542_ (
    .A(\memory[5][7] ),
    .B(_06147_),
    .Y(_00415_)
  );
  NAND _08543_ (
    .A(\memory[21][7] ),
    .B(_06167_),
    .Y(_00416_)
  );
  NAND _08544_ (
    .A(\memory[8][7] ),
    .B(_06374_),
    .Y(_00417_)
  );
  NAND _08545_ (
    .A(\memory[20][7] ),
    .B(_05930_),
    .Y(_00418_)
  );
  NAND _08546_ (
    .A(\memory[10][7] ),
    .B(_05899_),
    .Y(_00419_)
  );
  NAND _08547_ (
    .A(\memory[26][7] ),
    .B(_06333_),
    .Y(_00420_)
  );
  NAND _08548_ (
    .A(\memory[4][7] ),
    .B(_05961_),
    .Y(_00421_)
  );
  NAND _08549_ (
    .A(\memory[16][7] ),
    .B(_06085_),
    .Y(_00422_)
  );
  NAND _08550_ (
    .A(\memory[28][7] ),
    .B(_05981_),
    .Y(_00423_)
  );
  AND _08551_ (
    .A(_00400_),
    .B(_00409_),
    .Y(_00424_)
  );
  AND _08552_ (
    .A(_00404_),
    .B(_00420_),
    .Y(_00425_)
  );
  AND _08553_ (
    .A(_00396_),
    .B(_00402_),
    .Y(_00426_)
  );
  AND _08554_ (
    .A(_00418_),
    .B(_00422_),
    .Y(_00427_)
  );
  AND _08555_ (
    .A(_00426_),
    .B(_00427_),
    .Y(_00428_)
  );
  AND _08556_ (
    .A(_00414_),
    .B(_00424_),
    .Y(_00429_)
  );
  AND _08557_ (
    .A(_00411_),
    .B(_00429_),
    .Y(_00430_)
  );
  AND _08558_ (
    .A(_00428_),
    .B(_00430_),
    .Y(_00431_)
  );
  AND _08559_ (
    .A(_00398_),
    .B(_00401_),
    .Y(_00432_)
  );
  AND _08560_ (
    .A(_00397_),
    .B(_00432_),
    .Y(_00433_)
  );
  AND _08561_ (
    .A(_00425_),
    .B(_00433_),
    .Y(_00434_)
  );
  AND _08562_ (
    .A(_00392_),
    .B(_00415_),
    .Y(_00435_)
  );
  AND _08563_ (
    .A(_00399_),
    .B(_00417_),
    .Y(_00436_)
  );
  AND _08564_ (
    .A(_00435_),
    .B(_00436_),
    .Y(_00437_)
  );
  AND _08565_ (
    .A(_00434_),
    .B(_00437_),
    .Y(_00438_)
  );
  AND _08566_ (
    .A(_00431_),
    .B(_00438_),
    .Y(_00439_)
  );
  AND _08567_ (
    .A(_00393_),
    .B(_00419_),
    .Y(_00440_)
  );
  AND _08568_ (
    .A(_00391_),
    .B(_00416_),
    .Y(_00441_)
  );
  AND _08569_ (
    .A(_00423_),
    .B(_00441_),
    .Y(_00442_)
  );
  AND _08570_ (
    .A(_00440_),
    .B(_00442_),
    .Y(_00443_)
  );
  AND _08571_ (
    .A(_00412_),
    .B(_00443_),
    .Y(_00444_)
  );
  AND _08572_ (
    .A(_00403_),
    .B(_00405_),
    .Y(_00445_)
  );
  AND _08573_ (
    .A(_00394_),
    .B(_00445_),
    .Y(_00446_)
  );
  AND _08574_ (
    .A(_00395_),
    .B(_00413_),
    .Y(_00447_)
  );
  AND _08575_ (
    .A(_00410_),
    .B(_00447_),
    .Y(_00448_)
  );
  AND _08576_ (
    .A(_00408_),
    .B(_00421_),
    .Y(_00449_)
  );
  AND _08577_ (
    .A(_00448_),
    .B(_00449_),
    .Y(_00450_)
  );
  AND _08578_ (
    .A(_00446_),
    .B(_00450_),
    .Y(_00451_)
  );
  AND _08579_ (
    .A(_00444_),
    .B(_00451_),
    .Y(_00452_)
  );
  NAND _08580_ (
    .A(_00439_),
    .B(_00452_),
    .Y(\data_mem_o[23] )
  );
  NAND _08581_ (
    .A(\memory[29][0] ),
    .B(_05826_),
    .Y(_00453_)
  );
  NAND _08582_ (
    .A(\memory[13][0] ),
    .B(_06002_),
    .Y(_00454_)
  );
  NAND _08583_ (
    .A(\memory[14][0] ),
    .B(_06064_),
    .Y(_00455_)
  );
  AND _08584_ (
    .A(_00454_),
    .B(_00455_),
    .Y(_00456_)
  );
  AND _08585_ (
    .A(_00453_),
    .B(_00456_),
    .Y(_00457_)
  );
  NAND _08586_ (
    .A(\memory[2][0] ),
    .B(_05599_),
    .Y(_00458_)
  );
  NAND _08587_ (
    .A(\memory[18][0] ),
    .B(_05754_),
    .Y(_00459_)
  );
  AND _08588_ (
    .A(_00458_),
    .B(_00459_),
    .Y(_00460_)
  );
  NAND _08589_ (
    .A(\memory[28][0] ),
    .B(_05847_),
    .Y(_00461_)
  );
  NAND _08590_ (
    .A(\memory[30][0] ),
    .B(_05692_),
    .Y(_00462_)
  );
  AND _08591_ (
    .A(_00461_),
    .B(_00462_),
    .Y(_00463_)
  );
  AND _08592_ (
    .A(_00460_),
    .B(_00463_),
    .Y(_00464_)
  );
  NAND _08593_ (
    .A(\memory[1][0] ),
    .B(_06043_),
    .Y(_00465_)
  );
  NAND _08594_ (
    .A(\memory[17][0] ),
    .B(_05558_),
    .Y(_00466_)
  );
  AND _08595_ (
    .A(_00465_),
    .B(_00466_),
    .Y(_00467_)
  );
  NAND _08596_ (
    .A(\memory[6][0] ),
    .B(_05475_),
    .Y(_00468_)
  );
  NAND _08597_ (
    .A(\memory[21][0] ),
    .B(_05806_),
    .Y(_00469_)
  );
  AND _08598_ (
    .A(_00468_),
    .B(_00469_),
    .Y(_00470_)
  );
  AND _08599_ (
    .A(_00467_),
    .B(_00470_),
    .Y(_00471_)
  );
  AND _08600_ (
    .A(_00464_),
    .B(_00471_),
    .Y(_00472_)
  );
  AND _08601_ (
    .A(_00457_),
    .B(_00472_),
    .Y(_00473_)
  );
  NAND _08602_ (
    .A(\memory[27][0] ),
    .B(_05981_),
    .Y(_00474_)
  );
  NAND _08603_ (
    .A(\memory[15][0] ),
    .B(_06085_),
    .Y(_00475_)
  );
  AND _08604_ (
    .A(_00474_),
    .B(_00475_),
    .Y(_00476_)
  );
  NAND _08605_ (
    .A(\memory[25][0] ),
    .B(_06333_),
    .Y(_00477_)
  );
  NAND _08606_ (
    .A(\memory[7][0] ),
    .B(_06374_),
    .Y(_00478_)
  );
  AND _08607_ (
    .A(_00477_),
    .B(_00478_),
    .Y(_00479_)
  );
  AND _08608_ (
    .A(_00476_),
    .B(_00479_),
    .Y(_00480_)
  );
  NAND _08609_ (
    .A(\memory[5][0] ),
    .B(_05733_),
    .Y(_00481_)
  );
  NAND _08610_ (
    .A(\memory[11][0] ),
    .B(_05661_),
    .Y(_00482_)
  );
  AND _08611_ (
    .A(_00481_),
    .B(_00482_),
    .Y(_00483_)
  );
  NAND _08612_ (
    .A(\memory[12][0] ),
    .B(_05785_),
    .Y(_00484_)
  );
  NAND _08613_ (
    .A(\memory[22][0] ),
    .B(_06023_),
    .Y(_00485_)
  );
  AND _08614_ (
    .A(_00484_),
    .B(_00485_),
    .Y(_00486_)
  );
  AND _08615_ (
    .A(_00483_),
    .B(_00486_),
    .Y(_00487_)
  );
  NAND _08616_ (
    .A(\memory[10][0] ),
    .B(_06312_),
    .Y(_00488_)
  );
  NAND _08617_ (
    .A(\memory[31][0] ),
    .B(_06188_),
    .Y(_00489_)
  );
  NAND _08618_ (
    .A(\memory[16][0] ),
    .B(_06209_),
    .Y(_00490_)
  );
  AND _08619_ (
    .A(_00489_),
    .B(_00490_),
    .Y(_00491_)
  );
  NAND _08620_ (
    .A(\memory[0][0] ),
    .B(_06116_),
    .Y(_00492_)
  );
  NAND _08621_ (
    .A(\memory[20][0] ),
    .B(_06167_),
    .Y(_00493_)
  );
  NAND _08622_ (
    .A(\memory[4][0] ),
    .B(_06147_),
    .Y(_00494_)
  );
  AND _08623_ (
    .A(_00493_),
    .B(_00494_),
    .Y(_00495_)
  );
  AND _08624_ (
    .A(_00492_),
    .B(_00495_),
    .Y(_00496_)
  );
  AND _08625_ (
    .A(_00491_),
    .B(_00496_),
    .Y(_00497_)
  );
  AND _08626_ (
    .A(_00488_),
    .B(_00497_),
    .Y(_00498_)
  );
  AND _08627_ (
    .A(_00487_),
    .B(_00498_),
    .Y(_00499_)
  );
  AND _08628_ (
    .A(_00480_),
    .B(_00499_),
    .Y(_00500_)
  );
  NAND _08629_ (
    .A(\memory[19][0] ),
    .B(_05930_),
    .Y(_00501_)
  );
  NAND _08630_ (
    .A(\memory[26][0] ),
    .B(_06291_),
    .Y(_00502_)
  );
  NAND _08631_ (
    .A(\memory[24][0] ),
    .B(_06250_),
    .Y(_00503_)
  );
  AND _08632_ (
    .A(_00502_),
    .B(_00503_),
    .Y(_00504_)
  );
  AND _08633_ (
    .A(_00501_),
    .B(_00504_),
    .Y(_00505_)
  );
  NAND _08634_ (
    .A(\memory[8][0] ),
    .B(_06353_),
    .Y(_00506_)
  );
  NAND _08635_ (
    .A(\memory[9][0] ),
    .B(_05899_),
    .Y(_00507_)
  );
  AND _08636_ (
    .A(_00506_),
    .B(_00507_),
    .Y(_00508_)
  );
  NAND _08637_ (
    .A(\memory[3][0] ),
    .B(_05961_),
    .Y(_00509_)
  );
  NAND _08638_ (
    .A(\memory[23][0] ),
    .B(_06395_),
    .Y(_00510_)
  );
  AND _08639_ (
    .A(_00509_),
    .B(_00510_),
    .Y(_00511_)
  );
  AND _08640_ (
    .A(_00508_),
    .B(_00511_),
    .Y(_00512_)
  );
  AND _08641_ (
    .A(_00505_),
    .B(_00512_),
    .Y(_00513_)
  );
  AND _08642_ (
    .A(_00500_),
    .B(_00513_),
    .Y(_00514_)
  );
  NAND _08643_ (
    .A(_00473_),
    .B(_00514_),
    .Y(\data_mem_o[8] )
  );
  NAND _08644_ (
    .A(\memory[5][1] ),
    .B(_05733_),
    .Y(_00515_)
  );
  NAND _08645_ (
    .A(\memory[2][1] ),
    .B(_05599_),
    .Y(_00516_)
  );
  NAND _08646_ (
    .A(\memory[18][1] ),
    .B(_05754_),
    .Y(_00517_)
  );
  NAND _08647_ (
    .A(\memory[29][1] ),
    .B(_05826_),
    .Y(_00518_)
  );
  NAND _08648_ (
    .A(\memory[14][1] ),
    .B(_06064_),
    .Y(_00519_)
  );
  NAND _08649_ (
    .A(\memory[21][1] ),
    .B(_05806_),
    .Y(_00520_)
  );
  NAND _08650_ (
    .A(\memory[6][1] ),
    .B(_05475_),
    .Y(_00521_)
  );
  NAND _08651_ (
    .A(\memory[28][1] ),
    .B(_05847_),
    .Y(_00522_)
  );
  NAND _08652_ (
    .A(\memory[11][1] ),
    .B(_05661_),
    .Y(_00523_)
  );
  NAND _08653_ (
    .A(\memory[30][1] ),
    .B(_05692_),
    .Y(_00524_)
  );
  NAND _08654_ (
    .A(\memory[1][1] ),
    .B(_06043_),
    .Y(_00525_)
  );
  NAND _08655_ (
    .A(\memory[23][1] ),
    .B(_06395_),
    .Y(_00526_)
  );
  NAND _08656_ (
    .A(\memory[24][1] ),
    .B(_06250_),
    .Y(_00527_)
  );
  NAND _08657_ (
    .A(\memory[26][1] ),
    .B(_06291_),
    .Y(_00528_)
  );
  NAND _08658_ (
    .A(\memory[27][1] ),
    .B(_05981_),
    .Y(_00529_)
  );
  NAND _08659_ (
    .A(\memory[17][1] ),
    .B(_05558_),
    .Y(_00530_)
  );
  NAND _08660_ (
    .A(\memory[13][1] ),
    .B(_06002_),
    .Y(_00531_)
  );
  NAND _08661_ (
    .A(\memory[22][1] ),
    .B(_06023_),
    .Y(_00532_)
  );
  NAND _08662_ (
    .A(\memory[12][1] ),
    .B(_05785_),
    .Y(_00533_)
  );
  NAND _08663_ (
    .A(\memory[9][1] ),
    .B(_05899_),
    .Y(_00534_)
  );
  NAND _08664_ (
    .A(\memory[16][1] ),
    .B(_06209_),
    .Y(_00535_)
  );
  NAND _08665_ (
    .A(\memory[20][1] ),
    .B(_06167_),
    .Y(_00536_)
  );
  NAND _08666_ (
    .A(\memory[4][1] ),
    .B(_06147_),
    .Y(_00537_)
  );
  NAND _08667_ (
    .A(\memory[31][1] ),
    .B(_06188_),
    .Y(_00538_)
  );
  NAND _08668_ (
    .A(\memory[0][1] ),
    .B(_06116_),
    .Y(_00539_)
  );
  NAND _08669_ (
    .A(\memory[8][1] ),
    .B(_06353_),
    .Y(_00540_)
  );
  NAND _08670_ (
    .A(\memory[19][1] ),
    .B(_05930_),
    .Y(_00541_)
  );
  NAND _08671_ (
    .A(\memory[7][1] ),
    .B(_06374_),
    .Y(_00542_)
  );
  NAND _08672_ (
    .A(\memory[25][1] ),
    .B(_06333_),
    .Y(_00543_)
  );
  NAND _08673_ (
    .A(\memory[15][1] ),
    .B(_06085_),
    .Y(_00544_)
  );
  NAND _08674_ (
    .A(\memory[3][1] ),
    .B(_05961_),
    .Y(_00545_)
  );
  NAND _08675_ (
    .A(\memory[10][1] ),
    .B(_06312_),
    .Y(_00546_)
  );
  AND _08676_ (
    .A(_00519_),
    .B(_00531_),
    .Y(_00547_)
  );
  AND _08677_ (
    .A(_00522_),
    .B(_00524_),
    .Y(_00548_)
  );
  AND _08678_ (
    .A(_00520_),
    .B(_00532_),
    .Y(_00549_)
  );
  AND _08679_ (
    .A(_00521_),
    .B(_00526_),
    .Y(_00550_)
  );
  AND _08680_ (
    .A(_00549_),
    .B(_00550_),
    .Y(_00551_)
  );
  AND _08681_ (
    .A(_00516_),
    .B(_00540_),
    .Y(_00552_)
  );
  AND _08682_ (
    .A(_00518_),
    .B(_00536_),
    .Y(_00553_)
  );
  AND _08683_ (
    .A(_00515_),
    .B(_00553_),
    .Y(_00554_)
  );
  AND _08684_ (
    .A(_00552_),
    .B(_00554_),
    .Y(_00555_)
  );
  AND _08685_ (
    .A(_00551_),
    .B(_00555_),
    .Y(_00556_)
  );
  AND _08686_ (
    .A(_00535_),
    .B(_00556_),
    .Y(_00557_)
  );
  AND _08687_ (
    .A(_00528_),
    .B(_00543_),
    .Y(_00558_)
  );
  AND _08688_ (
    .A(_00527_),
    .B(_00548_),
    .Y(_00559_)
  );
  AND _08689_ (
    .A(_00558_),
    .B(_00559_),
    .Y(_00560_)
  );
  AND _08690_ (
    .A(_00529_),
    .B(_00530_),
    .Y(_00561_)
  );
  AND _08691_ (
    .A(_00538_),
    .B(_00561_),
    .Y(_00562_)
  );
  AND _08692_ (
    .A(_00517_),
    .B(_00541_),
    .Y(_00563_)
  );
  AND _08693_ (
    .A(_00539_),
    .B(_00563_),
    .Y(_00564_)
  );
  AND _08694_ (
    .A(_00562_),
    .B(_00564_),
    .Y(_00565_)
  );
  AND _08695_ (
    .A(_00560_),
    .B(_00565_),
    .Y(_00566_)
  );
  AND _08696_ (
    .A(_00542_),
    .B(_00545_),
    .Y(_00567_)
  );
  AND _08697_ (
    .A(_00525_),
    .B(_00567_),
    .Y(_00568_)
  );
  AND _08698_ (
    .A(_00523_),
    .B(_00533_),
    .Y(_00569_)
  );
  AND _08699_ (
    .A(_00537_),
    .B(_00569_),
    .Y(_00570_)
  );
  AND _08700_ (
    .A(_00547_),
    .B(_00570_),
    .Y(_00571_)
  );
  AND _08701_ (
    .A(_00534_),
    .B(_00544_),
    .Y(_00572_)
  );
  AND _08702_ (
    .A(_00546_),
    .B(_00572_),
    .Y(_00573_)
  );
  AND _08703_ (
    .A(_00571_),
    .B(_00573_),
    .Y(_00574_)
  );
  AND _08704_ (
    .A(_00568_),
    .B(_00574_),
    .Y(_00575_)
  );
  AND _08705_ (
    .A(_00566_),
    .B(_00575_),
    .Y(_00576_)
  );
  NAND _08706_ (
    .A(_00557_),
    .B(_00576_),
    .Y(\data_mem_o[9] )
  );
  NAND _08707_ (
    .A(\memory[22][2] ),
    .B(_06023_),
    .Y(_00577_)
  );
  NAND _08708_ (
    .A(\memory[21][2] ),
    .B(_05806_),
    .Y(_00578_)
  );
  NAND _08709_ (
    .A(\memory[29][2] ),
    .B(_05826_),
    .Y(_00579_)
  );
  NAND _08710_ (
    .A(\memory[18][2] ),
    .B(_05754_),
    .Y(_00580_)
  );
  NAND _08711_ (
    .A(\memory[2][2] ),
    .B(_05599_),
    .Y(_00581_)
  );
  NAND _08712_ (
    .A(\memory[1][2] ),
    .B(_06043_),
    .Y(_00582_)
  );
  NAND _08713_ (
    .A(\memory[12][2] ),
    .B(_05785_),
    .Y(_00583_)
  );
  NAND _08714_ (
    .A(\memory[28][2] ),
    .B(_05847_),
    .Y(_00584_)
  );
  NAND _08715_ (
    .A(\memory[14][2] ),
    .B(_06064_),
    .Y(_00585_)
  );
  NAND _08716_ (
    .A(\memory[30][2] ),
    .B(_05692_),
    .Y(_00586_)
  );
  NAND _08717_ (
    .A(\memory[13][2] ),
    .B(_06002_),
    .Y(_00587_)
  );
  NAND _08718_ (
    .A(\memory[24][2] ),
    .B(_06250_),
    .Y(_00588_)
  );
  NAND _08719_ (
    .A(\memory[15][2] ),
    .B(_06085_),
    .Y(_00589_)
  );
  NAND _08720_ (
    .A(\memory[25][2] ),
    .B(_06333_),
    .Y(_00590_)
  );
  NAND _08721_ (
    .A(\memory[3][2] ),
    .B(_05961_),
    .Y(_00591_)
  );
  NAND _08722_ (
    .A(\memory[5][2] ),
    .B(_05733_),
    .Y(_00592_)
  );
  NAND _08723_ (
    .A(\memory[11][2] ),
    .B(_05661_),
    .Y(_00593_)
  );
  NAND _08724_ (
    .A(\memory[17][2] ),
    .B(_05558_),
    .Y(_00594_)
  );
  NAND _08725_ (
    .A(\memory[6][2] ),
    .B(_05475_),
    .Y(_00595_)
  );
  NAND _08726_ (
    .A(\memory[7][2] ),
    .B(_06374_),
    .Y(_00596_)
  );
  NAND _08727_ (
    .A(\memory[0][2] ),
    .B(_06116_),
    .Y(_00597_)
  );
  NAND _08728_ (
    .A(\memory[20][2] ),
    .B(_06167_),
    .Y(_00598_)
  );
  NAND _08729_ (
    .A(\memory[4][2] ),
    .B(_06147_),
    .Y(_00599_)
  );
  NAND _08730_ (
    .A(\memory[16][2] ),
    .B(_06209_),
    .Y(_00600_)
  );
  NAND _08731_ (
    .A(\memory[31][2] ),
    .B(_06188_),
    .Y(_00601_)
  );
  NAND _08732_ (
    .A(\memory[9][2] ),
    .B(_05899_),
    .Y(_00602_)
  );
  NAND _08733_ (
    .A(\memory[10][2] ),
    .B(_06312_),
    .Y(_00603_)
  );
  NAND _08734_ (
    .A(\memory[26][2] ),
    .B(_06291_),
    .Y(_00604_)
  );
  NAND _08735_ (
    .A(\memory[27][2] ),
    .B(_05981_),
    .Y(_00605_)
  );
  NAND _08736_ (
    .A(\memory[19][2] ),
    .B(_05930_),
    .Y(_00606_)
  );
  NAND _08737_ (
    .A(\memory[23][2] ),
    .B(_06395_),
    .Y(_00607_)
  );
  NAND _08738_ (
    .A(\memory[8][2] ),
    .B(_06353_),
    .Y(_00608_)
  );
  AND _08739_ (
    .A(_00584_),
    .B(_00586_),
    .Y(_00609_)
  );
  AND _08740_ (
    .A(_00577_),
    .B(_00578_),
    .Y(_00610_)
  );
  AND _08741_ (
    .A(_00600_),
    .B(_00607_),
    .Y(_00611_)
  );
  AND _08742_ (
    .A(_00610_),
    .B(_00611_),
    .Y(_00612_)
  );
  AND _08743_ (
    .A(_00602_),
    .B(_00603_),
    .Y(_00613_)
  );
  AND _08744_ (
    .A(_00579_),
    .B(_00598_),
    .Y(_00614_)
  );
  AND _08745_ (
    .A(_00583_),
    .B(_00614_),
    .Y(_00615_)
  );
  AND _08746_ (
    .A(_00613_),
    .B(_00615_),
    .Y(_00616_)
  );
  AND _08747_ (
    .A(_00612_),
    .B(_00616_),
    .Y(_00617_)
  );
  AND _08748_ (
    .A(_00582_),
    .B(_00617_),
    .Y(_00618_)
  );
  AND _08749_ (
    .A(_00590_),
    .B(_00604_),
    .Y(_00619_)
  );
  AND _08750_ (
    .A(_00588_),
    .B(_00609_),
    .Y(_00620_)
  );
  AND _08751_ (
    .A(_00619_),
    .B(_00620_),
    .Y(_00621_)
  );
  AND _08752_ (
    .A(_00594_),
    .B(_00605_),
    .Y(_00622_)
  );
  AND _08753_ (
    .A(_00601_),
    .B(_00622_),
    .Y(_00623_)
  );
  AND _08754_ (
    .A(_00580_),
    .B(_00606_),
    .Y(_00624_)
  );
  AND _08755_ (
    .A(_00597_),
    .B(_00624_),
    .Y(_00625_)
  );
  AND _08756_ (
    .A(_00623_),
    .B(_00625_),
    .Y(_00626_)
  );
  AND _08757_ (
    .A(_00621_),
    .B(_00626_),
    .Y(_00627_)
  );
  AND _08758_ (
    .A(_00581_),
    .B(_00591_),
    .Y(_00628_)
  );
  AND _08759_ (
    .A(_00592_),
    .B(_00599_),
    .Y(_00629_)
  );
  AND _08760_ (
    .A(_00596_),
    .B(_00629_),
    .Y(_00630_)
  );
  AND _08761_ (
    .A(_00595_),
    .B(_00630_),
    .Y(_00631_)
  );
  AND _08762_ (
    .A(_00587_),
    .B(_00593_),
    .Y(_00632_)
  );
  AND _08763_ (
    .A(_00589_),
    .B(_00632_),
    .Y(_00633_)
  );
  AND _08764_ (
    .A(_00585_),
    .B(_00608_),
    .Y(_00634_)
  );
  AND _08765_ (
    .A(_00633_),
    .B(_00634_),
    .Y(_00635_)
  );
  AND _08766_ (
    .A(_00631_),
    .B(_00635_),
    .Y(_00636_)
  );
  AND _08767_ (
    .A(_00628_),
    .B(_00636_),
    .Y(_00637_)
  );
  AND _08768_ (
    .A(_00627_),
    .B(_00637_),
    .Y(_00638_)
  );
  NAND _08769_ (
    .A(_00618_),
    .B(_00638_),
    .Y(\data_mem_o[10] )
  );
  NAND _08770_ (
    .A(\memory[13][3] ),
    .B(_06002_),
    .Y(_00639_)
  );
  NAND _08771_ (
    .A(\memory[1][3] ),
    .B(_06043_),
    .Y(_00640_)
  );
  NAND _08772_ (
    .A(\memory[18][3] ),
    .B(_05754_),
    .Y(_00641_)
  );
  NAND _08773_ (
    .A(\memory[17][3] ),
    .B(_05558_),
    .Y(_00642_)
  );
  NAND _08774_ (
    .A(\memory[21][3] ),
    .B(_05806_),
    .Y(_00643_)
  );
  AND _08775_ (
    .A(_00642_),
    .B(_00643_),
    .Y(_00644_)
  );
  NAND _08776_ (
    .A(\memory[30][3] ),
    .B(_05692_),
    .Y(_00645_)
  );
  NAND _08777_ (
    .A(\memory[2][3] ),
    .B(_05599_),
    .Y(_00646_)
  );
  NAND _08778_ (
    .A(\memory[11][3] ),
    .B(_05661_),
    .Y(_00647_)
  );
  NAND _08779_ (
    .A(\memory[29][3] ),
    .B(_05826_),
    .Y(_00648_)
  );
  NAND _08780_ (
    .A(\memory[14][3] ),
    .B(_06064_),
    .Y(_00649_)
  );
  NAND _08781_ (
    .A(\memory[6][3] ),
    .B(_05475_),
    .Y(_00650_)
  );
  NAND _08782_ (
    .A(\memory[15][3] ),
    .B(_06085_),
    .Y(_00651_)
  );
  NAND _08783_ (
    .A(\memory[25][3] ),
    .B(_06333_),
    .Y(_00652_)
  );
  AND _08784_ (
    .A(_00651_),
    .B(_00652_),
    .Y(_00653_)
  );
  NAND _08785_ (
    .A(\memory[3][3] ),
    .B(_05961_),
    .Y(_00654_)
  );
  NAND _08786_ (
    .A(\memory[26][3] ),
    .B(_06291_),
    .Y(_00655_)
  );
  NAND _08787_ (
    .A(\memory[28][3] ),
    .B(_05847_),
    .Y(_00656_)
  );
  NAND _08788_ (
    .A(\memory[22][3] ),
    .B(_06023_),
    .Y(_00657_)
  );
  NAND _08789_ (
    .A(\memory[12][3] ),
    .B(_05785_),
    .Y(_00658_)
  );
  NAND _08790_ (
    .A(\memory[5][3] ),
    .B(_05733_),
    .Y(_00659_)
  );
  NAND _08791_ (
    .A(\memory[9][3] ),
    .B(_05899_),
    .Y(_00660_)
  );
  NAND _08792_ (
    .A(\memory[0][3] ),
    .B(_06116_),
    .Y(_00661_)
  );
  NAND _08793_ (
    .A(\memory[4][3] ),
    .B(_06147_),
    .Y(_00662_)
  );
  NAND _08794_ (
    .A(\memory[20][3] ),
    .B(_06167_),
    .Y(_00663_)
  );
  NAND _08795_ (
    .A(\memory[16][3] ),
    .B(_06209_),
    .Y(_00664_)
  );
  NAND _08796_ (
    .A(\memory[31][3] ),
    .B(_06188_),
    .Y(_00665_)
  );
  NAND _08797_ (
    .A(\memory[7][3] ),
    .B(_06374_),
    .Y(_00666_)
  );
  NAND _08798_ (
    .A(\memory[24][3] ),
    .B(_06250_),
    .Y(_00667_)
  );
  NAND _08799_ (
    .A(\memory[8][3] ),
    .B(_06353_),
    .Y(_00668_)
  );
  NAND _08800_ (
    .A(\memory[27][3] ),
    .B(_05981_),
    .Y(_00669_)
  );
  NAND _08801_ (
    .A(\memory[19][3] ),
    .B(_05930_),
    .Y(_00670_)
  );
  AND _08802_ (
    .A(_00669_),
    .B(_00670_),
    .Y(_00671_)
  );
  NAND _08803_ (
    .A(\memory[10][3] ),
    .B(_06312_),
    .Y(_00672_)
  );
  NAND _08804_ (
    .A(\memory[23][3] ),
    .B(_06395_),
    .Y(_00673_)
  );
  AND _08805_ (
    .A(_00650_),
    .B(_00657_),
    .Y(_00674_)
  );
  AND _08806_ (
    .A(_00648_),
    .B(_00674_),
    .Y(_00675_)
  );
  AND _08807_ (
    .A(_00659_),
    .B(_00675_),
    .Y(_00676_)
  );
  AND _08808_ (
    .A(_00647_),
    .B(_00649_),
    .Y(_00677_)
  );
  AND _08809_ (
    .A(_00658_),
    .B(_00677_),
    .Y(_00678_)
  );
  AND _08810_ (
    .A(_00640_),
    .B(_00656_),
    .Y(_00679_)
  );
  AND _08811_ (
    .A(_00678_),
    .B(_00679_),
    .Y(_00680_)
  );
  AND _08812_ (
    .A(_00676_),
    .B(_00680_),
    .Y(_00681_)
  );
  AND _08813_ (
    .A(_00661_),
    .B(_00664_),
    .Y(_00682_)
  );
  AND _08814_ (
    .A(_00639_),
    .B(_00682_),
    .Y(_00683_)
  );
  AND _08815_ (
    .A(_00663_),
    .B(_00665_),
    .Y(_00684_)
  );
  AND _08816_ (
    .A(_00662_),
    .B(_00684_),
    .Y(_00685_)
  );
  AND _08817_ (
    .A(_00683_),
    .B(_00685_),
    .Y(_00686_)
  );
  AND _08818_ (
    .A(_00653_),
    .B(_00686_),
    .Y(_00687_)
  );
  AND _08819_ (
    .A(_00641_),
    .B(_00673_),
    .Y(_00688_)
  );
  AND _08820_ (
    .A(_00671_),
    .B(_00688_),
    .Y(_00689_)
  );
  AND _08821_ (
    .A(_00687_),
    .B(_00689_),
    .Y(_00690_)
  );
  AND _08822_ (
    .A(_00681_),
    .B(_00690_),
    .Y(_00691_)
  );
  AND _08823_ (
    .A(_00644_),
    .B(_00645_),
    .Y(_00692_)
  );
  AND _08824_ (
    .A(_00660_),
    .B(_00672_),
    .Y(_00693_)
  );
  AND _08825_ (
    .A(_00654_),
    .B(_00666_),
    .Y(_00694_)
  );
  AND _08826_ (
    .A(_00693_),
    .B(_00694_),
    .Y(_00695_)
  );
  AND _08827_ (
    .A(_00646_),
    .B(_00668_),
    .Y(_00696_)
  );
  AND _08828_ (
    .A(_00655_),
    .B(_00667_),
    .Y(_00697_)
  );
  AND _08829_ (
    .A(_00696_),
    .B(_00697_),
    .Y(_00698_)
  );
  AND _08830_ (
    .A(_00695_),
    .B(_00698_),
    .Y(_00699_)
  );
  AND _08831_ (
    .A(_00692_),
    .B(_00699_),
    .Y(_00700_)
  );
  NAND _08832_ (
    .A(_00691_),
    .B(_00700_),
    .Y(\data_mem_o[11] )
  );
  NAND _08833_ (
    .A(\memory[22][4] ),
    .B(_06023_),
    .Y(_00701_)
  );
  NAND _08834_ (
    .A(\memory[21][4] ),
    .B(_05806_),
    .Y(_00702_)
  );
  NAND _08835_ (
    .A(\memory[2][4] ),
    .B(_05599_),
    .Y(_00703_)
  );
  NAND _08836_ (
    .A(\memory[28][4] ),
    .B(_05847_),
    .Y(_00704_)
  );
  NAND _08837_ (
    .A(\memory[30][4] ),
    .B(_05692_),
    .Y(_00705_)
  );
  NAND _08838_ (
    .A(\memory[29][4] ),
    .B(_05826_),
    .Y(_00706_)
  );
  NAND _08839_ (
    .A(\memory[18][4] ),
    .B(_05754_),
    .Y(_00707_)
  );
  NAND _08840_ (
    .A(\memory[6][4] ),
    .B(_05475_),
    .Y(_00708_)
  );
  NAND _08841_ (
    .A(\memory[13][4] ),
    .B(_06002_),
    .Y(_00709_)
  );
  NAND _08842_ (
    .A(\memory[5][4] ),
    .B(_05733_),
    .Y(_00710_)
  );
  NAND _08843_ (
    .A(\memory[17][4] ),
    .B(_05558_),
    .Y(_00711_)
  );
  NAND _08844_ (
    .A(\memory[27][4] ),
    .B(_05981_),
    .Y(_00712_)
  );
  NAND _08845_ (
    .A(\memory[23][4] ),
    .B(_06395_),
    .Y(_00713_)
  );
  NAND _08846_ (
    .A(\memory[15][4] ),
    .B(_06085_),
    .Y(_00714_)
  );
  NAND _08847_ (
    .A(\memory[19][4] ),
    .B(_05930_),
    .Y(_00715_)
  );
  NAND _08848_ (
    .A(\memory[12][4] ),
    .B(_05785_),
    .Y(_00716_)
  );
  NAND _08849_ (
    .A(\memory[14][4] ),
    .B(_06064_),
    .Y(_00717_)
  );
  NAND _08850_ (
    .A(\memory[11][4] ),
    .B(_05661_),
    .Y(_00718_)
  );
  NAND _08851_ (
    .A(\memory[1][4] ),
    .B(_06043_),
    .Y(_00719_)
  );
  NAND _08852_ (
    .A(\memory[10][4] ),
    .B(_06312_),
    .Y(_00720_)
  );
  NAND _08853_ (
    .A(\memory[16][4] ),
    .B(_06209_),
    .Y(_00721_)
  );
  NAND _08854_ (
    .A(\memory[20][4] ),
    .B(_06167_),
    .Y(_00722_)
  );
  NAND _08855_ (
    .A(\memory[4][4] ),
    .B(_06147_),
    .Y(_00723_)
  );
  NAND _08856_ (
    .A(\memory[31][4] ),
    .B(_06188_),
    .Y(_00724_)
  );
  NAND _08857_ (
    .A(\memory[0][4] ),
    .B(_06116_),
    .Y(_00725_)
  );
  NAND _08858_ (
    .A(\memory[24][4] ),
    .B(_06250_),
    .Y(_00726_)
  );
  NAND _08859_ (
    .A(\memory[9][4] ),
    .B(_05899_),
    .Y(_00727_)
  );
  NAND _08860_ (
    .A(\memory[7][4] ),
    .B(_06374_),
    .Y(_00728_)
  );
  NAND _08861_ (
    .A(\memory[26][4] ),
    .B(_06291_),
    .Y(_00729_)
  );
  NAND _08862_ (
    .A(\memory[8][4] ),
    .B(_06353_),
    .Y(_00730_)
  );
  NAND _08863_ (
    .A(\memory[25][4] ),
    .B(_06333_),
    .Y(_00731_)
  );
  NAND _08864_ (
    .A(\memory[3][4] ),
    .B(_05961_),
    .Y(_00732_)
  );
  AND _08865_ (
    .A(_00701_),
    .B(_00702_),
    .Y(_00733_)
  );
  AND _08866_ (
    .A(_00731_),
    .B(_00733_),
    .Y(_00734_)
  );
  AND _08867_ (
    .A(_00706_),
    .B(_00722_),
    .Y(_00735_)
  );
  AND _08868_ (
    .A(_00729_),
    .B(_00735_),
    .Y(_00736_)
  );
  AND _08869_ (
    .A(_00734_),
    .B(_00736_),
    .Y(_00737_)
  );
  AND _08870_ (
    .A(_00714_),
    .B(_00718_),
    .Y(_00738_)
  );
  AND _08871_ (
    .A(_00720_),
    .B(_00727_),
    .Y(_00739_)
  );
  AND _08872_ (
    .A(_00738_),
    .B(_00739_),
    .Y(_00740_)
  );
  AND _08873_ (
    .A(_00737_),
    .B(_00740_),
    .Y(_00741_)
  );
  AND _08874_ (
    .A(_00710_),
    .B(_00723_),
    .Y(_00742_)
  );
  AND _08875_ (
    .A(_00728_),
    .B(_00742_),
    .Y(_00743_)
  );
  AND _08876_ (
    .A(_00708_),
    .B(_00743_),
    .Y(_00744_)
  );
  AND _08877_ (
    .A(_00709_),
    .B(_00717_),
    .Y(_00745_)
  );
  AND _08878_ (
    .A(_00716_),
    .B(_00745_),
    .Y(_00746_)
  );
  AND _08879_ (
    .A(_00721_),
    .B(_00746_),
    .Y(_00747_)
  );
  AND _08880_ (
    .A(_00744_),
    .B(_00747_),
    .Y(_00748_)
  );
  AND _08881_ (
    .A(_00741_),
    .B(_00748_),
    .Y(_00749_)
  );
  AND _08882_ (
    .A(_00711_),
    .B(_00712_),
    .Y(_00750_)
  );
  AND _08883_ (
    .A(_00724_),
    .B(_00750_),
    .Y(_00751_)
  );
  AND _08884_ (
    .A(_00704_),
    .B(_00715_),
    .Y(_00752_)
  );
  AND _08885_ (
    .A(_00725_),
    .B(_00752_),
    .Y(_00753_)
  );
  AND _08886_ (
    .A(_00751_),
    .B(_00753_),
    .Y(_00754_)
  );
  AND _08887_ (
    .A(_00705_),
    .B(_00707_),
    .Y(_00755_)
  );
  AND _08888_ (
    .A(_00713_),
    .B(_00726_),
    .Y(_00756_)
  );
  AND _08889_ (
    .A(_00755_),
    .B(_00756_),
    .Y(_00757_)
  );
  AND _08890_ (
    .A(_00703_),
    .B(_00732_),
    .Y(_00758_)
  );
  AND _08891_ (
    .A(_00719_),
    .B(_00730_),
    .Y(_00759_)
  );
  AND _08892_ (
    .A(_00758_),
    .B(_00759_),
    .Y(_00760_)
  );
  AND _08893_ (
    .A(_00757_),
    .B(_00760_),
    .Y(_00761_)
  );
  AND _08894_ (
    .A(_00754_),
    .B(_00761_),
    .Y(_00762_)
  );
  NAND _08895_ (
    .A(_00749_),
    .B(_00762_),
    .Y(\data_mem_o[12] )
  );
  NAND _08896_ (
    .A(\memory[12][5] ),
    .B(_05785_),
    .Y(_00763_)
  );
  NAND _08897_ (
    .A(\memory[11][5] ),
    .B(_05661_),
    .Y(_00764_)
  );
  NAND _08898_ (
    .A(\memory[18][5] ),
    .B(_05754_),
    .Y(_00765_)
  );
  NAND _08899_ (
    .A(\memory[2][5] ),
    .B(_05599_),
    .Y(_00766_)
  );
  NAND _08900_ (
    .A(\memory[13][5] ),
    .B(_06002_),
    .Y(_00767_)
  );
  NAND _08901_ (
    .A(\memory[1][5] ),
    .B(_06043_),
    .Y(_00768_)
  );
  NAND _08902_ (
    .A(\memory[30][5] ),
    .B(_05692_),
    .Y(_00769_)
  );
  NAND _08903_ (
    .A(\memory[5][5] ),
    .B(_05733_),
    .Y(_00770_)
  );
  NAND _08904_ (
    .A(\memory[29][5] ),
    .B(_05826_),
    .Y(_00771_)
  );
  NAND _08905_ (
    .A(\memory[14][5] ),
    .B(_06064_),
    .Y(_00772_)
  );
  NAND _08906_ (
    .A(\memory[28][5] ),
    .B(_05847_),
    .Y(_00773_)
  );
  NAND _08907_ (
    .A(\memory[8][5] ),
    .B(_06353_),
    .Y(_00774_)
  );
  NAND _08908_ (
    .A(\memory[15][5] ),
    .B(_06085_),
    .Y(_00775_)
  );
  NAND _08909_ (
    .A(\memory[9][5] ),
    .B(_05899_),
    .Y(_00776_)
  );
  NAND _08910_ (
    .A(\memory[3][5] ),
    .B(_05961_),
    .Y(_00777_)
  );
  NAND _08911_ (
    .A(\memory[17][5] ),
    .B(_05558_),
    .Y(_00778_)
  );
  NAND _08912_ (
    .A(\memory[6][5] ),
    .B(_05475_),
    .Y(_00779_)
  );
  NAND _08913_ (
    .A(\memory[22][5] ),
    .B(_06023_),
    .Y(_00780_)
  );
  NAND _08914_ (
    .A(\memory[21][5] ),
    .B(_05806_),
    .Y(_00781_)
  );
  NAND _08915_ (
    .A(\memory[27][5] ),
    .B(_05981_),
    .Y(_00782_)
  );
  NAND _08916_ (
    .A(\memory[31][5] ),
    .B(_06188_),
    .Y(_00783_)
  );
  NAND _08917_ (
    .A(\memory[16][5] ),
    .B(_06209_),
    .Y(_00784_)
  );
  NAND _08918_ (
    .A(\memory[0][5] ),
    .B(_06116_),
    .Y(_00785_)
  );
  NAND _08919_ (
    .A(\memory[20][5] ),
    .B(_06167_),
    .Y(_00786_)
  );
  NAND _08920_ (
    .A(\memory[4][5] ),
    .B(_06147_),
    .Y(_00787_)
  );
  NAND _08921_ (
    .A(\memory[25][5] ),
    .B(_06333_),
    .Y(_00788_)
  );
  NAND _08922_ (
    .A(\memory[19][5] ),
    .B(_05930_),
    .Y(_00789_)
  );
  NAND _08923_ (
    .A(\memory[24][5] ),
    .B(_06250_),
    .Y(_00790_)
  );
  NAND _08924_ (
    .A(\memory[7][5] ),
    .B(_06374_),
    .Y(_00791_)
  );
  NAND _08925_ (
    .A(\memory[23][5] ),
    .B(_06395_),
    .Y(_00792_)
  );
  NAND _08926_ (
    .A(\memory[10][5] ),
    .B(_06312_),
    .Y(_00793_)
  );
  NAND _08927_ (
    .A(\memory[26][5] ),
    .B(_06291_),
    .Y(_00794_)
  );
  AND _08928_ (
    .A(_00767_),
    .B(_00780_),
    .Y(_00795_)
  );
  AND _08929_ (
    .A(_00772_),
    .B(_00781_),
    .Y(_00796_)
  );
  AND _08930_ (
    .A(_00795_),
    .B(_00796_),
    .Y(_00797_)
  );
  AND _08931_ (
    .A(_00765_),
    .B(_00790_),
    .Y(_00798_)
  );
  AND _08932_ (
    .A(_00768_),
    .B(_00774_),
    .Y(_00799_)
  );
  AND _08933_ (
    .A(_00786_),
    .B(_00791_),
    .Y(_00800_)
  );
  AND _08934_ (
    .A(_00788_),
    .B(_00800_),
    .Y(_00801_)
  );
  AND _08935_ (
    .A(_00770_),
    .B(_00787_),
    .Y(_00802_)
  );
  AND _08936_ (
    .A(_00782_),
    .B(_00802_),
    .Y(_00803_)
  );
  AND _08937_ (
    .A(_00801_),
    .B(_00803_),
    .Y(_00804_)
  );
  AND _08938_ (
    .A(_00799_),
    .B(_00804_),
    .Y(_00805_)
  );
  AND _08939_ (
    .A(_00764_),
    .B(_00776_),
    .Y(_00806_)
  );
  AND _08940_ (
    .A(_00783_),
    .B(_00806_),
    .Y(_00807_)
  );
  AND _08941_ (
    .A(_00769_),
    .B(_00785_),
    .Y(_00808_)
  );
  AND _08942_ (
    .A(_00766_),
    .B(_00777_),
    .Y(_00809_)
  );
  AND _08943_ (
    .A(_00808_),
    .B(_00809_),
    .Y(_00810_)
  );
  AND _08944_ (
    .A(_00807_),
    .B(_00810_),
    .Y(_00811_)
  );
  AND _08945_ (
    .A(_00789_),
    .B(_00798_),
    .Y(_00812_)
  );
  AND _08946_ (
    .A(_00763_),
    .B(_00784_),
    .Y(_00813_)
  );
  AND _08947_ (
    .A(_00793_),
    .B(_00813_),
    .Y(_00814_)
  );
  AND _08948_ (
    .A(_00812_),
    .B(_00814_),
    .Y(_00815_)
  );
  AND _08949_ (
    .A(_00811_),
    .B(_00815_),
    .Y(_00816_)
  );
  AND _08950_ (
    .A(_00778_),
    .B(_00792_),
    .Y(_00817_)
  );
  AND _08951_ (
    .A(_00775_),
    .B(_00779_),
    .Y(_00818_)
  );
  AND _08952_ (
    .A(_00817_),
    .B(_00818_),
    .Y(_00819_)
  );
  AND _08953_ (
    .A(_00797_),
    .B(_00819_),
    .Y(_00820_)
  );
  AND _08954_ (
    .A(_00771_),
    .B(_00794_),
    .Y(_00821_)
  );
  AND _08955_ (
    .A(_00773_),
    .B(_00821_),
    .Y(_00822_)
  );
  AND _08956_ (
    .A(_00820_),
    .B(_00822_),
    .Y(_00823_)
  );
  AND _08957_ (
    .A(_00816_),
    .B(_00823_),
    .Y(_00824_)
  );
  NAND _08958_ (
    .A(_00805_),
    .B(_00824_),
    .Y(\data_mem_o[13] )
  );
  NAND _08959_ (
    .A(\memory[11][6] ),
    .B(_05661_),
    .Y(_00825_)
  );
  NAND _08960_ (
    .A(\memory[6][6] ),
    .B(_05475_),
    .Y(_00826_)
  );
  NAND _08961_ (
    .A(\memory[18][6] ),
    .B(_05754_),
    .Y(_00827_)
  );
  NAND _08962_ (
    .A(\memory[1][6] ),
    .B(_06043_),
    .Y(_00828_)
  );
  NAND _08963_ (
    .A(\memory[5][6] ),
    .B(_05733_),
    .Y(_00829_)
  );
  AND _08964_ (
    .A(_00828_),
    .B(_00829_),
    .Y(_00830_)
  );
  NAND _08965_ (
    .A(\memory[30][6] ),
    .B(_05692_),
    .Y(_00831_)
  );
  NAND _08966_ (
    .A(\memory[29][6] ),
    .B(_05826_),
    .Y(_00832_)
  );
  NAND _08967_ (
    .A(\memory[12][6] ),
    .B(_05785_),
    .Y(_00833_)
  );
  NAND _08968_ (
    .A(\memory[13][6] ),
    .B(_06002_),
    .Y(_00834_)
  );
  NAND _08969_ (
    .A(\memory[2][6] ),
    .B(_05599_),
    .Y(_00835_)
  );
  NAND _08970_ (
    .A(\memory[14][6] ),
    .B(_06064_),
    .Y(_00836_)
  );
  NAND _08971_ (
    .A(\memory[8][6] ),
    .B(_06353_),
    .Y(_00837_)
  );
  NAND _08972_ (
    .A(\memory[9][6] ),
    .B(_05899_),
    .Y(_00838_)
  );
  NAND _08973_ (
    .A(\memory[27][6] ),
    .B(_05981_),
    .Y(_00839_)
  );
  NAND _08974_ (
    .A(\memory[3][6] ),
    .B(_05961_),
    .Y(_00840_)
  );
  NAND _08975_ (
    .A(\memory[21][6] ),
    .B(_05806_),
    .Y(_00841_)
  );
  NAND _08976_ (
    .A(\memory[17][6] ),
    .B(_05558_),
    .Y(_00842_)
  );
  AND _08977_ (
    .A(_00841_),
    .B(_00842_),
    .Y(_00843_)
  );
  NAND _08978_ (
    .A(\memory[22][6] ),
    .B(_06023_),
    .Y(_00844_)
  );
  NAND _08979_ (
    .A(\memory[28][6] ),
    .B(_05847_),
    .Y(_00845_)
  );
  NAND _08980_ (
    .A(\memory[15][6] ),
    .B(_06085_),
    .Y(_00846_)
  );
  NAND _08981_ (
    .A(\memory[31][6] ),
    .B(_06188_),
    .Y(_00847_)
  );
  NAND _08982_ (
    .A(\memory[20][6] ),
    .B(_06167_),
    .Y(_00848_)
  );
  NAND _08983_ (
    .A(\memory[4][6] ),
    .B(_06147_),
    .Y(_00849_)
  );
  NAND _08984_ (
    .A(\memory[0][6] ),
    .B(_06116_),
    .Y(_00850_)
  );
  NAND _08985_ (
    .A(\memory[16][6] ),
    .B(_06209_),
    .Y(_00851_)
  );
  NAND _08986_ (
    .A(\memory[7][6] ),
    .B(_06374_),
    .Y(_00852_)
  );
  NAND _08987_ (
    .A(\memory[19][6] ),
    .B(_05930_),
    .Y(_00853_)
  );
  NAND _08988_ (
    .A(\memory[26][6] ),
    .B(_06291_),
    .Y(_00854_)
  );
  NAND _08989_ (
    .A(\memory[25][6] ),
    .B(_06333_),
    .Y(_00855_)
  );
  NAND _08990_ (
    .A(\memory[23][6] ),
    .B(_06395_),
    .Y(_00856_)
  );
  NAND _08991_ (
    .A(\memory[24][6] ),
    .B(_06250_),
    .Y(_00857_)
  );
  NAND _08992_ (
    .A(\memory[10][6] ),
    .B(_06312_),
    .Y(_00858_)
  );
  AND _08993_ (
    .A(_00832_),
    .B(_00843_),
    .Y(_00859_)
  );
  AND _08994_ (
    .A(_00845_),
    .B(_00859_),
    .Y(_00860_)
  );
  AND _08995_ (
    .A(_00834_),
    .B(_00836_),
    .Y(_00861_)
  );
  AND _08996_ (
    .A(_00833_),
    .B(_00844_),
    .Y(_00862_)
  );
  AND _08997_ (
    .A(_00861_),
    .B(_00862_),
    .Y(_00863_)
  );
  AND _08998_ (
    .A(_00860_),
    .B(_00863_),
    .Y(_00864_)
  );
  AND _08999_ (
    .A(_00848_),
    .B(_00850_),
    .Y(_00865_)
  );
  AND _09000_ (
    .A(_00826_),
    .B(_00865_),
    .Y(_00866_)
  );
  AND _09001_ (
    .A(_00847_),
    .B(_00851_),
    .Y(_00867_)
  );
  AND _09002_ (
    .A(_00849_),
    .B(_00867_),
    .Y(_00868_)
  );
  AND _09003_ (
    .A(_00866_),
    .B(_00868_),
    .Y(_00869_)
  );
  AND _09004_ (
    .A(_00835_),
    .B(_00838_),
    .Y(_00870_)
  );
  AND _09005_ (
    .A(_00869_),
    .B(_00870_),
    .Y(_00871_)
  );
  AND _09006_ (
    .A(_00827_),
    .B(_00857_),
    .Y(_00872_)
  );
  AND _09007_ (
    .A(_00856_),
    .B(_00858_),
    .Y(_00873_)
  );
  AND _09008_ (
    .A(_00872_),
    .B(_00873_),
    .Y(_00874_)
  );
  AND _09009_ (
    .A(_00871_),
    .B(_00874_),
    .Y(_00875_)
  );
  AND _09010_ (
    .A(_00864_),
    .B(_00875_),
    .Y(_00876_)
  );
  AND _09011_ (
    .A(_00825_),
    .B(_00830_),
    .Y(_00877_)
  );
  AND _09012_ (
    .A(_00831_),
    .B(_00877_),
    .Y(_00878_)
  );
  AND _09013_ (
    .A(_00837_),
    .B(_00855_),
    .Y(_00879_)
  );
  AND _09014_ (
    .A(_00839_),
    .B(_00852_),
    .Y(_00880_)
  );
  AND _09015_ (
    .A(_00879_),
    .B(_00880_),
    .Y(_00881_)
  );
  AND _09016_ (
    .A(_00840_),
    .B(_00853_),
    .Y(_00882_)
  );
  AND _09017_ (
    .A(_00846_),
    .B(_00854_),
    .Y(_00883_)
  );
  AND _09018_ (
    .A(_00882_),
    .B(_00883_),
    .Y(_00884_)
  );
  AND _09019_ (
    .A(_00881_),
    .B(_00884_),
    .Y(_00885_)
  );
  AND _09020_ (
    .A(_00878_),
    .B(_00885_),
    .Y(_00886_)
  );
  NAND _09021_ (
    .A(_00876_),
    .B(_00886_),
    .Y(\data_mem_o[14] )
  );
  NAND _09022_ (
    .A(\memory[22][7] ),
    .B(_06023_),
    .Y(_00887_)
  );
  NAND _09023_ (
    .A(\memory[18][7] ),
    .B(_05754_),
    .Y(_00888_)
  );
  NAND _09024_ (
    .A(\memory[17][7] ),
    .B(_05558_),
    .Y(_00889_)
  );
  NAND _09025_ (
    .A(\memory[11][7] ),
    .B(_05661_),
    .Y(_00890_)
  );
  NAND _09026_ (
    .A(\memory[1][7] ),
    .B(_06043_),
    .Y(_00891_)
  );
  NAND _09027_ (
    .A(\memory[28][7] ),
    .B(_05847_),
    .Y(_00892_)
  );
  NAND _09028_ (
    .A(\memory[29][7] ),
    .B(_05826_),
    .Y(_00893_)
  );
  NAND _09029_ (
    .A(\memory[12][7] ),
    .B(_05785_),
    .Y(_00894_)
  );
  NAND _09030_ (
    .A(\memory[21][7] ),
    .B(_05806_),
    .Y(_00895_)
  );
  NAND _09031_ (
    .A(\memory[5][7] ),
    .B(_05733_),
    .Y(_00896_)
  );
  NAND _09032_ (
    .A(\memory[6][7] ),
    .B(_05475_),
    .Y(_00897_)
  );
  NAND _09033_ (
    .A(\memory[8][7] ),
    .B(_06353_),
    .Y(_00898_)
  );
  NAND _09034_ (
    .A(\memory[3][7] ),
    .B(_05961_),
    .Y(_00899_)
  );
  NAND _09035_ (
    .A(\memory[24][7] ),
    .B(_06250_),
    .Y(_00900_)
  );
  NAND _09036_ (
    .A(\memory[19][7] ),
    .B(_05930_),
    .Y(_00901_)
  );
  NAND _09037_ (
    .A(\memory[13][7] ),
    .B(_06002_),
    .Y(_00902_)
  );
  NAND _09038_ (
    .A(\memory[2][7] ),
    .B(_05599_),
    .Y(_00903_)
  );
  NAND _09039_ (
    .A(\memory[14][7] ),
    .B(_06064_),
    .Y(_00904_)
  );
  NAND _09040_ (
    .A(\memory[30][7] ),
    .B(_05692_),
    .Y(_00905_)
  );
  NAND _09041_ (
    .A(\memory[15][7] ),
    .B(_06085_),
    .Y(_00906_)
  );
  NAND _09042_ (
    .A(\memory[0][7] ),
    .B(_06116_),
    .Y(_00907_)
  );
  NAND _09043_ (
    .A(\memory[20][7] ),
    .B(_06167_),
    .Y(_00908_)
  );
  NAND _09044_ (
    .A(\memory[4][7] ),
    .B(_06147_),
    .Y(_00909_)
  );
  NAND _09045_ (
    .A(\memory[16][7] ),
    .B(_06209_),
    .Y(_00910_)
  );
  NAND _09046_ (
    .A(\memory[31][7] ),
    .B(_06188_),
    .Y(_00911_)
  );
  NAND _09047_ (
    .A(\memory[10][7] ),
    .B(_06312_),
    .Y(_00912_)
  );
  NAND _09048_ (
    .A(\memory[9][7] ),
    .B(_05899_),
    .Y(_00913_)
  );
  AND _09049_ (
    .A(_00912_),
    .B(_00913_),
    .Y(_00914_)
  );
  NAND _09050_ (
    .A(\memory[7][7] ),
    .B(_06374_),
    .Y(_00915_)
  );
  NAND _09051_ (
    .A(\memory[25][7] ),
    .B(_06333_),
    .Y(_00916_)
  );
  NAND _09052_ (
    .A(\memory[26][7] ),
    .B(_06291_),
    .Y(_00917_)
  );
  NAND _09053_ (
    .A(\memory[23][7] ),
    .B(_06395_),
    .Y(_00918_)
  );
  NAND _09054_ (
    .A(\memory[27][7] ),
    .B(_05981_),
    .Y(_00919_)
  );
  AND _09055_ (
    .A(_00900_),
    .B(_00918_),
    .Y(_00920_)
  );
  AND _09056_ (
    .A(_00902_),
    .B(_00904_),
    .Y(_00921_)
  );
  AND _09057_ (
    .A(_00894_),
    .B(_00921_),
    .Y(_00922_)
  );
  AND _09058_ (
    .A(_00910_),
    .B(_00922_),
    .Y(_00923_)
  );
  AND _09059_ (
    .A(_00898_),
    .B(_00923_),
    .Y(_00924_)
  );
  AND _09060_ (
    .A(_00888_),
    .B(_00905_),
    .Y(_00925_)
  );
  AND _09061_ (
    .A(_00920_),
    .B(_00925_),
    .Y(_00926_)
  );
  AND _09062_ (
    .A(_00889_),
    .B(_00919_),
    .Y(_00927_)
  );
  AND _09063_ (
    .A(_00911_),
    .B(_00927_),
    .Y(_00928_)
  );
  AND _09064_ (
    .A(_00892_),
    .B(_00901_),
    .Y(_00929_)
  );
  AND _09065_ (
    .A(_00907_),
    .B(_00929_),
    .Y(_00930_)
  );
  AND _09066_ (
    .A(_00928_),
    .B(_00930_),
    .Y(_00931_)
  );
  AND _09067_ (
    .A(_00926_),
    .B(_00931_),
    .Y(_00932_)
  );
  AND _09068_ (
    .A(_00887_),
    .B(_00895_),
    .Y(_00933_)
  );
  AND _09069_ (
    .A(_00916_),
    .B(_00933_),
    .Y(_00934_)
  );
  AND _09070_ (
    .A(_00893_),
    .B(_00908_),
    .Y(_00935_)
  );
  AND _09071_ (
    .A(_00917_),
    .B(_00935_),
    .Y(_00936_)
  );
  AND _09072_ (
    .A(_00934_),
    .B(_00936_),
    .Y(_00937_)
  );
  AND _09073_ (
    .A(_00890_),
    .B(_00906_),
    .Y(_00938_)
  );
  AND _09074_ (
    .A(_00914_),
    .B(_00938_),
    .Y(_00939_)
  );
  AND _09075_ (
    .A(_00937_),
    .B(_00939_),
    .Y(_00940_)
  );
  AND _09076_ (
    .A(_00899_),
    .B(_00903_),
    .Y(_00941_)
  );
  AND _09077_ (
    .A(_00896_),
    .B(_00909_),
    .Y(_00942_)
  );
  AND _09078_ (
    .A(_00915_),
    .B(_00942_),
    .Y(_00943_)
  );
  AND _09079_ (
    .A(_00891_),
    .B(_00897_),
    .Y(_00944_)
  );
  AND _09080_ (
    .A(_00943_),
    .B(_00944_),
    .Y(_00945_)
  );
  AND _09081_ (
    .A(_00941_),
    .B(_00945_),
    .Y(_00946_)
  );
  AND _09082_ (
    .A(_00940_),
    .B(_00946_),
    .Y(_00947_)
  );
  AND _09083_ (
    .A(_00932_),
    .B(_00947_),
    .Y(_00948_)
  );
  NAND _09084_ (
    .A(_00924_),
    .B(_00948_),
    .Y(\data_mem_o[15] )
  );
  NAND _09085_ (
    .A(\memory[21][0] ),
    .B(_06023_),
    .Y(_00949_)
  );
  NAND _09086_ (
    .A(\memory[17][0] ),
    .B(_05754_),
    .Y(_00950_)
  );
  NAND _09087_ (
    .A(\memory[12][0] ),
    .B(_06002_),
    .Y(_00951_)
  );
  NAND _09088_ (
    .A(\memory[20][0] ),
    .B(_05806_),
    .Y(_00952_)
  );
  NAND _09089_ (
    .A(\memory[28][0] ),
    .B(_05826_),
    .Y(_00953_)
  );
  NAND _09090_ (
    .A(\memory[1][0] ),
    .B(_05599_),
    .Y(_00954_)
  );
  NAND _09091_ (
    .A(\memory[4][0] ),
    .B(_05733_),
    .Y(_00955_)
  );
  NAND _09092_ (
    .A(\memory[11][0] ),
    .B(_05785_),
    .Y(_00956_)
  );
  NAND _09093_ (
    .A(\memory[29][0] ),
    .B(_05692_),
    .Y(_00957_)
  );
  NAND _09094_ (
    .A(\memory[10][0] ),
    .B(_05661_),
    .Y(_00958_)
  );
  NAND _09095_ (
    .A(\memory[27][0] ),
    .B(_05847_),
    .Y(_00959_)
  );
  NAND _09096_ (
    .A(\memory[8][0] ),
    .B(_05899_),
    .Y(_00960_)
  );
  NAND _09097_ (
    .A(\memory[26][0] ),
    .B(_05981_),
    .Y(_00961_)
  );
  NAND _09098_ (
    .A(\memory[6][0] ),
    .B(_06374_),
    .Y(_00962_)
  );
  NAND _09099_ (
    .A(\memory[18][0] ),
    .B(_05930_),
    .Y(_00963_)
  );
  NAND _09100_ (
    .A(\memory[13][0] ),
    .B(_06064_),
    .Y(_00964_)
  );
  NAND _09101_ (
    .A(\memory[16][0] ),
    .B(_05558_),
    .Y(_00965_)
  );
  NAND _09102_ (
    .A(\memory[5][0] ),
    .B(_05475_),
    .Y(_00966_)
  );
  NAND _09103_ (
    .A(\memory[0][0] ),
    .B(_06043_),
    .Y(_00967_)
  );
  NAND _09104_ (
    .A(\memory[9][0] ),
    .B(_06312_),
    .Y(_00968_)
  );
  NAND _09105_ (
    .A(\memory[30][0] ),
    .B(_06188_),
    .Y(_00969_)
  );
  NAND _09106_ (
    .A(\memory[15][0] ),
    .B(_06209_),
    .Y(_00970_)
  );
  NAND _09107_ (
    .A(\memory[31][0] ),
    .B(_06116_),
    .Y(_00971_)
  );
  NAND _09108_ (
    .A(\memory[3][0] ),
    .B(_06147_),
    .Y(_00972_)
  );
  NAND _09109_ (
    .A(\memory[19][0] ),
    .B(_06167_),
    .Y(_00973_)
  );
  NAND _09110_ (
    .A(\memory[22][0] ),
    .B(_06395_),
    .Y(_00974_)
  );
  NAND _09111_ (
    .A(\memory[14][0] ),
    .B(_06085_),
    .Y(_00975_)
  );
  NAND _09112_ (
    .A(\memory[23][0] ),
    .B(_06250_),
    .Y(_00976_)
  );
  NAND _09113_ (
    .A(\memory[2][0] ),
    .B(_05961_),
    .Y(_00977_)
  );
  NAND _09114_ (
    .A(\memory[7][0] ),
    .B(_06353_),
    .Y(_00978_)
  );
  NAND _09115_ (
    .A(\memory[24][0] ),
    .B(_06333_),
    .Y(_00979_)
  );
  NAND _09116_ (
    .A(\memory[25][0] ),
    .B(_06291_),
    .Y(_00980_)
  );
  AND _09117_ (
    .A(_00960_),
    .B(_00978_),
    .Y(_00981_)
  );
  AND _09118_ (
    .A(_00951_),
    .B(_00956_),
    .Y(_00982_)
  );
  AND _09119_ (
    .A(_00974_),
    .B(_00977_),
    .Y(_00983_)
  );
  AND _09120_ (
    .A(_00954_),
    .B(_00983_),
    .Y(_00984_)
  );
  AND _09121_ (
    .A(_00955_),
    .B(_00972_),
    .Y(_00985_)
  );
  AND _09122_ (
    .A(_00968_),
    .B(_00985_),
    .Y(_00986_)
  );
  AND _09123_ (
    .A(_00952_),
    .B(_00973_),
    .Y(_00987_)
  );
  AND _09124_ (
    .A(_00958_),
    .B(_00987_),
    .Y(_00988_)
  );
  AND _09125_ (
    .A(_00986_),
    .B(_00988_),
    .Y(_00989_)
  );
  AND _09126_ (
    .A(_00962_),
    .B(_00989_),
    .Y(_00990_)
  );
  AND _09127_ (
    .A(_00984_),
    .B(_00990_),
    .Y(_00991_)
  );
  AND _09128_ (
    .A(_00950_),
    .B(_00963_),
    .Y(_00992_)
  );
  AND _09129_ (
    .A(_00959_),
    .B(_00971_),
    .Y(_00993_)
  );
  AND _09130_ (
    .A(_00964_),
    .B(_00993_),
    .Y(_00994_)
  );
  AND _09131_ (
    .A(_00992_),
    .B(_00994_),
    .Y(_00995_)
  );
  AND _09132_ (
    .A(_00953_),
    .B(_00975_),
    .Y(_00996_)
  );
  AND _09133_ (
    .A(_00969_),
    .B(_00996_),
    .Y(_00997_)
  );
  AND _09134_ (
    .A(_00995_),
    .B(_00997_),
    .Y(_00998_)
  );
  AND _09135_ (
    .A(_00979_),
    .B(_00982_),
    .Y(_00999_)
  );
  AND _09136_ (
    .A(_00976_),
    .B(_00999_),
    .Y(_01000_)
  );
  AND _09137_ (
    .A(_00949_),
    .B(_01000_),
    .Y(_01001_)
  );
  AND _09138_ (
    .A(_00998_),
    .B(_01001_),
    .Y(_01002_)
  );
  AND _09139_ (
    .A(_00957_),
    .B(_00970_),
    .Y(_01003_)
  );
  AND _09140_ (
    .A(_00961_),
    .B(_01003_),
    .Y(_01004_)
  );
  AND _09141_ (
    .A(_00966_),
    .B(_01004_),
    .Y(_01005_)
  );
  AND _09142_ (
    .A(_00981_),
    .B(_01005_),
    .Y(_01006_)
  );
  AND _09143_ (
    .A(_00967_),
    .B(_00980_),
    .Y(_01007_)
  );
  AND _09144_ (
    .A(_00965_),
    .B(_01007_),
    .Y(_01008_)
  );
  AND _09145_ (
    .A(_01006_),
    .B(_01008_),
    .Y(_01009_)
  );
  AND _09146_ (
    .A(_01002_),
    .B(_01009_),
    .Y(_01010_)
  );
  NAND _09147_ (
    .A(_00991_),
    .B(_01010_),
    .Y(\data_mem_o[0] )
  );
  NAND _09148_ (
    .A(\memory[0][1] ),
    .B(_06043_),
    .Y(_01011_)
  );
  NAND _09149_ (
    .A(\memory[11][1] ),
    .B(_05785_),
    .Y(_01012_)
  );
  NAND _09150_ (
    .A(\memory[17][1] ),
    .B(_05754_),
    .Y(_01013_)
  );
  NAND _09151_ (
    .A(\memory[20][1] ),
    .B(_05806_),
    .Y(_01014_)
  );
  NAND _09152_ (
    .A(\memory[28][1] ),
    .B(_05826_),
    .Y(_01015_)
  );
  AND _09153_ (
    .A(_01014_),
    .B(_01015_),
    .Y(_01016_)
  );
  NAND _09154_ (
    .A(\memory[12][1] ),
    .B(_06002_),
    .Y(_01017_)
  );
  NAND _09155_ (
    .A(\memory[1][1] ),
    .B(_05599_),
    .Y(_01018_)
  );
  NAND _09156_ (
    .A(\memory[16][1] ),
    .B(_05558_),
    .Y(_01019_)
  );
  NAND _09157_ (
    .A(\memory[27][1] ),
    .B(_05847_),
    .Y(_01020_)
  );
  NAND _09158_ (
    .A(\memory[5][1] ),
    .B(_05475_),
    .Y(_01021_)
  );
  NAND _09159_ (
    .A(\memory[29][1] ),
    .B(_05692_),
    .Y(_01022_)
  );
  NAND _09160_ (
    .A(\memory[25][1] ),
    .B(_06291_),
    .Y(_01023_)
  );
  NAND _09161_ (
    .A(\memory[24][1] ),
    .B(_06333_),
    .Y(_01024_)
  );
  NAND _09162_ (
    .A(\memory[26][1] ),
    .B(_05981_),
    .Y(_01025_)
  );
  NAND _09163_ (
    .A(\memory[14][1] ),
    .B(_06085_),
    .Y(_01026_)
  );
  NAND _09164_ (
    .A(\memory[21][1] ),
    .B(_06023_),
    .Y(_01027_)
  );
  NAND _09165_ (
    .A(\memory[10][1] ),
    .B(_05661_),
    .Y(_01028_)
  );
  NAND _09166_ (
    .A(\memory[4][1] ),
    .B(_05733_),
    .Y(_01029_)
  );
  NAND _09167_ (
    .A(\memory[13][1] ),
    .B(_06064_),
    .Y(_01030_)
  );
  NAND _09168_ (
    .A(\memory[23][1] ),
    .B(_06250_),
    .Y(_01031_)
  );
  NAND _09169_ (
    .A(\memory[31][1] ),
    .B(_06116_),
    .Y(_01032_)
  );
  NAND _09170_ (
    .A(\memory[3][1] ),
    .B(_06147_),
    .Y(_01033_)
  );
  NAND _09171_ (
    .A(\memory[19][1] ),
    .B(_06167_),
    .Y(_01034_)
  );
  NAND _09172_ (
    .A(\memory[15][1] ),
    .B(_06209_),
    .Y(_01035_)
  );
  NAND _09173_ (
    .A(\memory[30][1] ),
    .B(_06188_),
    .Y(_01036_)
  );
  NAND _09174_ (
    .A(\memory[6][1] ),
    .B(_06374_),
    .Y(_01037_)
  );
  NAND _09175_ (
    .A(\memory[8][1] ),
    .B(_05899_),
    .Y(_01038_)
  );
  NAND _09176_ (
    .A(\memory[22][1] ),
    .B(_06395_),
    .Y(_01039_)
  );
  NAND _09177_ (
    .A(\memory[7][1] ),
    .B(_06353_),
    .Y(_01040_)
  );
  NAND _09178_ (
    .A(\memory[9][1] ),
    .B(_06312_),
    .Y(_01041_)
  );
  NAND _09179_ (
    .A(\memory[2][1] ),
    .B(_05961_),
    .Y(_01042_)
  );
  NAND _09180_ (
    .A(\memory[18][1] ),
    .B(_05930_),
    .Y(_01043_)
  );
  AND _09181_ (
    .A(_01041_),
    .B(_01042_),
    .Y(_01044_)
  );
  AND _09182_ (
    .A(_01011_),
    .B(_01012_),
    .Y(_01045_)
  );
  AND _09183_ (
    .A(_01017_),
    .B(_01045_),
    .Y(_01046_)
  );
  AND _09184_ (
    .A(_01021_),
    .B(_01025_),
    .Y(_01047_)
  );
  AND _09185_ (
    .A(_01037_),
    .B(_01040_),
    .Y(_01048_)
  );
  AND _09186_ (
    .A(_01035_),
    .B(_01048_),
    .Y(_01049_)
  );
  AND _09187_ (
    .A(_01047_),
    .B(_01049_),
    .Y(_01050_)
  );
  AND _09188_ (
    .A(_01031_),
    .B(_01046_),
    .Y(_01051_)
  );
  AND _09189_ (
    .A(_01016_),
    .B(_01023_),
    .Y(_01052_)
  );
  AND _09190_ (
    .A(_01051_),
    .B(_01052_),
    .Y(_01053_)
  );
  AND _09191_ (
    .A(_01050_),
    .B(_01053_),
    .Y(_01054_)
  );
  AND _09192_ (
    .A(_01018_),
    .B(_01027_),
    .Y(_01055_)
  );
  AND _09193_ (
    .A(_01024_),
    .B(_01055_),
    .Y(_01056_)
  );
  AND _09194_ (
    .A(_01019_),
    .B(_01038_),
    .Y(_01057_)
  );
  AND _09195_ (
    .A(_01028_),
    .B(_01057_),
    .Y(_01058_)
  );
  AND _09196_ (
    .A(_01056_),
    .B(_01058_),
    .Y(_01059_)
  );
  AND _09197_ (
    .A(_01013_),
    .B(_01036_),
    .Y(_01060_)
  );
  AND _09198_ (
    .A(_01059_),
    .B(_01060_),
    .Y(_01061_)
  );
  AND _09199_ (
    .A(_01054_),
    .B(_01061_),
    .Y(_01062_)
  );
  AND _09200_ (
    .A(_01032_),
    .B(_01033_),
    .Y(_01063_)
  );
  AND _09201_ (
    .A(_01039_),
    .B(_01063_),
    .Y(_01064_)
  );
  AND _09202_ (
    .A(_01029_),
    .B(_01064_),
    .Y(_01065_)
  );
  AND _09203_ (
    .A(_01022_),
    .B(_01026_),
    .Y(_01066_)
  );
  AND _09204_ (
    .A(_01020_),
    .B(_01034_),
    .Y(_01067_)
  );
  AND _09205_ (
    .A(_01030_),
    .B(_01067_),
    .Y(_01068_)
  );
  AND _09206_ (
    .A(_01066_),
    .B(_01068_),
    .Y(_01069_)
  );
  AND _09207_ (
    .A(_01043_),
    .B(_01069_),
    .Y(_01070_)
  );
  AND _09208_ (
    .A(_01044_),
    .B(_01070_),
    .Y(_01071_)
  );
  AND _09209_ (
    .A(_01065_),
    .B(_01071_),
    .Y(_01072_)
  );
  NAND _09210_ (
    .A(_01062_),
    .B(_01072_),
    .Y(\data_mem_o[1] )
  );
  NAND _09211_ (
    .A(\memory[0][2] ),
    .B(_06043_),
    .Y(_01073_)
  );
  NAND _09212_ (
    .A(\memory[11][2] ),
    .B(_05785_),
    .Y(_01074_)
  );
  NAND _09213_ (
    .A(\memory[17][2] ),
    .B(_05754_),
    .Y(_01075_)
  );
  AND _09214_ (
    .A(_01074_),
    .B(_01075_),
    .Y(_01076_)
  );
  AND _09215_ (
    .A(_01073_),
    .B(_01076_),
    .Y(_01077_)
  );
  NAND _09216_ (
    .A(\memory[20][2] ),
    .B(_05806_),
    .Y(_01078_)
  );
  NAND _09217_ (
    .A(\memory[28][2] ),
    .B(_05826_),
    .Y(_01079_)
  );
  AND _09218_ (
    .A(_01078_),
    .B(_01079_),
    .Y(_01080_)
  );
  NAND _09219_ (
    .A(\memory[12][2] ),
    .B(_06002_),
    .Y(_01081_)
  );
  NAND _09220_ (
    .A(\memory[1][2] ),
    .B(_05599_),
    .Y(_01082_)
  );
  AND _09221_ (
    .A(_01081_),
    .B(_01082_),
    .Y(_01083_)
  );
  AND _09222_ (
    .A(_01080_),
    .B(_01083_),
    .Y(_01084_)
  );
  NAND _09223_ (
    .A(\memory[16][2] ),
    .B(_05558_),
    .Y(_01085_)
  );
  NAND _09224_ (
    .A(\memory[27][2] ),
    .B(_05847_),
    .Y(_01086_)
  );
  AND _09225_ (
    .A(_01085_),
    .B(_01086_),
    .Y(_01087_)
  );
  NAND _09226_ (
    .A(\memory[5][2] ),
    .B(_05475_),
    .Y(_01088_)
  );
  NAND _09227_ (
    .A(\memory[29][2] ),
    .B(_05692_),
    .Y(_01089_)
  );
  AND _09228_ (
    .A(_01088_),
    .B(_01089_),
    .Y(_01090_)
  );
  AND _09229_ (
    .A(_01087_),
    .B(_01090_),
    .Y(_01091_)
  );
  AND _09230_ (
    .A(_01084_),
    .B(_01091_),
    .Y(_01092_)
  );
  AND _09231_ (
    .A(_01077_),
    .B(_01092_),
    .Y(_01093_)
  );
  NAND _09232_ (
    .A(\memory[25][2] ),
    .B(_06291_),
    .Y(_01094_)
  );
  NAND _09233_ (
    .A(\memory[24][2] ),
    .B(_06333_),
    .Y(_01095_)
  );
  AND _09234_ (
    .A(_01094_),
    .B(_01095_),
    .Y(_01096_)
  );
  NAND _09235_ (
    .A(\memory[26][2] ),
    .B(_05981_),
    .Y(_01097_)
  );
  NAND _09236_ (
    .A(\memory[9][2] ),
    .B(_06312_),
    .Y(_01098_)
  );
  AND _09237_ (
    .A(_01097_),
    .B(_01098_),
    .Y(_01099_)
  );
  AND _09238_ (
    .A(_01096_),
    .B(_01099_),
    .Y(_01100_)
  );
  NAND _09239_ (
    .A(\memory[21][2] ),
    .B(_06023_),
    .Y(_01101_)
  );
  NAND _09240_ (
    .A(\memory[10][2] ),
    .B(_05661_),
    .Y(_01102_)
  );
  AND _09241_ (
    .A(_01101_),
    .B(_01102_),
    .Y(_01103_)
  );
  NAND _09242_ (
    .A(\memory[13][2] ),
    .B(_06064_),
    .Y(_01104_)
  );
  NAND _09243_ (
    .A(\memory[4][2] ),
    .B(_05733_),
    .Y(_01105_)
  );
  AND _09244_ (
    .A(_01104_),
    .B(_01105_),
    .Y(_01106_)
  );
  AND _09245_ (
    .A(_01103_),
    .B(_01106_),
    .Y(_01107_)
  );
  NAND _09246_ (
    .A(\memory[23][2] ),
    .B(_06250_),
    .Y(_01108_)
  );
  NAND _09247_ (
    .A(\memory[31][2] ),
    .B(_06116_),
    .Y(_01109_)
  );
  NAND _09248_ (
    .A(\memory[3][2] ),
    .B(_06147_),
    .Y(_01110_)
  );
  NAND _09249_ (
    .A(\memory[19][2] ),
    .B(_06167_),
    .Y(_01111_)
  );
  AND _09250_ (
    .A(_01110_),
    .B(_01111_),
    .Y(_01112_)
  );
  AND _09251_ (
    .A(_01109_),
    .B(_01112_),
    .Y(_01113_)
  );
  NAND _09252_ (
    .A(\memory[15][2] ),
    .B(_06209_),
    .Y(_01114_)
  );
  NAND _09253_ (
    .A(\memory[30][2] ),
    .B(_06188_),
    .Y(_01115_)
  );
  AND _09254_ (
    .A(_01114_),
    .B(_01115_),
    .Y(_01116_)
  );
  AND _09255_ (
    .A(_01113_),
    .B(_01116_),
    .Y(_01117_)
  );
  AND _09256_ (
    .A(_01108_),
    .B(_01117_),
    .Y(_01118_)
  );
  AND _09257_ (
    .A(_01107_),
    .B(_01118_),
    .Y(_01119_)
  );
  AND _09258_ (
    .A(_01100_),
    .B(_01119_),
    .Y(_01120_)
  );
  NAND _09259_ (
    .A(\memory[14][2] ),
    .B(_06085_),
    .Y(_01121_)
  );
  NAND _09260_ (
    .A(\memory[6][2] ),
    .B(_06374_),
    .Y(_01122_)
  );
  NAND _09261_ (
    .A(\memory[22][2] ),
    .B(_06395_),
    .Y(_01123_)
  );
  AND _09262_ (
    .A(_01122_),
    .B(_01123_),
    .Y(_01124_)
  );
  AND _09263_ (
    .A(_01121_),
    .B(_01124_),
    .Y(_01125_)
  );
  NAND _09264_ (
    .A(\memory[8][2] ),
    .B(_05899_),
    .Y(_01126_)
  );
  NAND _09265_ (
    .A(\memory[18][2] ),
    .B(_05930_),
    .Y(_01127_)
  );
  AND _09266_ (
    .A(_01126_),
    .B(_01127_),
    .Y(_01128_)
  );
  NAND _09267_ (
    .A(\memory[7][2] ),
    .B(_06353_),
    .Y(_01129_)
  );
  NAND _09268_ (
    .A(\memory[2][2] ),
    .B(_05961_),
    .Y(_01130_)
  );
  AND _09269_ (
    .A(_01129_),
    .B(_01130_),
    .Y(_01131_)
  );
  AND _09270_ (
    .A(_01128_),
    .B(_01131_),
    .Y(_01132_)
  );
  AND _09271_ (
    .A(_01125_),
    .B(_01132_),
    .Y(_01133_)
  );
  AND _09272_ (
    .A(_01120_),
    .B(_01133_),
    .Y(_01134_)
  );
  NAND _09273_ (
    .A(_01093_),
    .B(_01134_),
    .Y(\data_mem_o[2] )
  );
  NAND _09274_ (
    .A(\memory[0][3] ),
    .B(_06043_),
    .Y(_01135_)
  );
  NAND _09275_ (
    .A(\memory[4][3] ),
    .B(_05733_),
    .Y(_01136_)
  );
  NAND _09276_ (
    .A(\memory[17][3] ),
    .B(_05754_),
    .Y(_01137_)
  );
  NAND _09277_ (
    .A(\memory[1][3] ),
    .B(_05599_),
    .Y(_01138_)
  );
  NAND _09278_ (
    .A(\memory[20][3] ),
    .B(_05806_),
    .Y(_01139_)
  );
  NAND _09279_ (
    .A(\memory[5][3] ),
    .B(_05475_),
    .Y(_01140_)
  );
  NAND _09280_ (
    .A(\memory[29][3] ),
    .B(_05692_),
    .Y(_01141_)
  );
  NAND _09281_ (
    .A(\memory[16][3] ),
    .B(_05558_),
    .Y(_01142_)
  );
  NAND _09282_ (
    .A(\memory[28][3] ),
    .B(_05826_),
    .Y(_01143_)
  );
  NAND _09283_ (
    .A(\memory[10][3] ),
    .B(_05661_),
    .Y(_01144_)
  );
  NAND _09284_ (
    .A(\memory[27][3] ),
    .B(_05847_),
    .Y(_01145_)
  );
  NAND _09285_ (
    .A(\memory[22][3] ),
    .B(_06395_),
    .Y(_01146_)
  );
  NAND _09286_ (
    .A(\memory[2][3] ),
    .B(_05961_),
    .Y(_01147_)
  );
  AND _09287_ (
    .A(_01146_),
    .B(_01147_),
    .Y(_01148_)
  );
  NAND _09288_ (
    .A(\memory[7][3] ),
    .B(_06353_),
    .Y(_01149_)
  );
  NAND _09289_ (
    .A(\memory[23][3] ),
    .B(_06250_),
    .Y(_01150_)
  );
  NAND _09290_ (
    .A(\memory[13][3] ),
    .B(_06064_),
    .Y(_01151_)
  );
  NAND _09291_ (
    .A(\memory[12][3] ),
    .B(_06002_),
    .Y(_01152_)
  );
  NAND _09292_ (
    .A(\memory[21][3] ),
    .B(_06023_),
    .Y(_01153_)
  );
  NAND _09293_ (
    .A(\memory[11][3] ),
    .B(_05785_),
    .Y(_01154_)
  );
  NAND _09294_ (
    .A(\memory[25][3] ),
    .B(_06291_),
    .Y(_01155_)
  );
  NAND _09295_ (
    .A(\memory[31][3] ),
    .B(_06116_),
    .Y(_01156_)
  );
  NAND _09296_ (
    .A(\memory[3][3] ),
    .B(_06147_),
    .Y(_01157_)
  );
  NAND _09297_ (
    .A(\memory[19][3] ),
    .B(_06167_),
    .Y(_01158_)
  );
  NAND _09298_ (
    .A(\memory[15][3] ),
    .B(_06209_),
    .Y(_01159_)
  );
  NAND _09299_ (
    .A(\memory[30][3] ),
    .B(_06188_),
    .Y(_01160_)
  );
  NAND _09300_ (
    .A(\memory[8][3] ),
    .B(_05899_),
    .Y(_01161_)
  );
  NAND _09301_ (
    .A(\memory[6][3] ),
    .B(_06374_),
    .Y(_01162_)
  );
  NAND _09302_ (
    .A(\memory[9][3] ),
    .B(_06312_),
    .Y(_01163_)
  );
  NAND _09303_ (
    .A(\memory[26][3] ),
    .B(_05981_),
    .Y(_01164_)
  );
  NAND _09304_ (
    .A(\memory[14][3] ),
    .B(_06085_),
    .Y(_01165_)
  );
  NAND _09305_ (
    .A(\memory[18][3] ),
    .B(_05930_),
    .Y(_01166_)
  );
  NAND _09306_ (
    .A(\memory[24][3] ),
    .B(_06333_),
    .Y(_01167_)
  );
  AND _09307_ (
    .A(_01152_),
    .B(_01154_),
    .Y(_01168_)
  );
  AND _09308_ (
    .A(_01149_),
    .B(_01161_),
    .Y(_01169_)
  );
  AND _09309_ (
    .A(_01141_),
    .B(_01159_),
    .Y(_01170_)
  );
  AND _09310_ (
    .A(_01164_),
    .B(_01170_),
    .Y(_01171_)
  );
  AND _09311_ (
    .A(_01140_),
    .B(_01171_),
    .Y(_01172_)
  );
  AND _09312_ (
    .A(_01169_),
    .B(_01172_),
    .Y(_01173_)
  );
  AND _09313_ (
    .A(_01135_),
    .B(_01155_),
    .Y(_01174_)
  );
  AND _09314_ (
    .A(_01142_),
    .B(_01174_),
    .Y(_01175_)
  );
  AND _09315_ (
    .A(_01173_),
    .B(_01175_),
    .Y(_01176_)
  );
  AND _09316_ (
    .A(_01138_),
    .B(_01148_),
    .Y(_01177_)
  );
  AND _09317_ (
    .A(_01136_),
    .B(_01157_),
    .Y(_01178_)
  );
  AND _09318_ (
    .A(_01163_),
    .B(_01178_),
    .Y(_01179_)
  );
  AND _09319_ (
    .A(_01139_),
    .B(_01158_),
    .Y(_01180_)
  );
  AND _09320_ (
    .A(_01144_),
    .B(_01180_),
    .Y(_01181_)
  );
  AND _09321_ (
    .A(_01179_),
    .B(_01181_),
    .Y(_01182_)
  );
  AND _09322_ (
    .A(_01162_),
    .B(_01182_),
    .Y(_01183_)
  );
  AND _09323_ (
    .A(_01177_),
    .B(_01183_),
    .Y(_01184_)
  );
  AND _09324_ (
    .A(_01176_),
    .B(_01184_),
    .Y(_01185_)
  );
  AND _09325_ (
    .A(_01137_),
    .B(_01166_),
    .Y(_01186_)
  );
  AND _09326_ (
    .A(_01145_),
    .B(_01156_),
    .Y(_01187_)
  );
  AND _09327_ (
    .A(_01151_),
    .B(_01187_),
    .Y(_01188_)
  );
  AND _09328_ (
    .A(_01186_),
    .B(_01188_),
    .Y(_01189_)
  );
  AND _09329_ (
    .A(_01143_),
    .B(_01165_),
    .Y(_01190_)
  );
  AND _09330_ (
    .A(_01160_),
    .B(_01190_),
    .Y(_01191_)
  );
  AND _09331_ (
    .A(_01167_),
    .B(_01168_),
    .Y(_01192_)
  );
  AND _09332_ (
    .A(_01150_),
    .B(_01192_),
    .Y(_01193_)
  );
  AND _09333_ (
    .A(_01153_),
    .B(_01193_),
    .Y(_01194_)
  );
  AND _09334_ (
    .A(_01191_),
    .B(_01194_),
    .Y(_01195_)
  );
  AND _09335_ (
    .A(_01189_),
    .B(_01195_),
    .Y(_01196_)
  );
  NAND _09336_ (
    .A(_01185_),
    .B(_01196_),
    .Y(\data_mem_o[3] )
  );
  NAND _09337_ (
    .A(\memory[21][4] ),
    .B(_06023_),
    .Y(_01197_)
  );
  NAND _09338_ (
    .A(\memory[17][4] ),
    .B(_05754_),
    .Y(_01198_)
  );
  NAND _09339_ (
    .A(\memory[12][4] ),
    .B(_06002_),
    .Y(_01199_)
  );
  NAND _09340_ (
    .A(\memory[20][4] ),
    .B(_05806_),
    .Y(_01200_)
  );
  NAND _09341_ (
    .A(\memory[28][4] ),
    .B(_05826_),
    .Y(_01201_)
  );
  NAND _09342_ (
    .A(\memory[1][4] ),
    .B(_05599_),
    .Y(_01202_)
  );
  NAND _09343_ (
    .A(\memory[4][4] ),
    .B(_05733_),
    .Y(_01203_)
  );
  NAND _09344_ (
    .A(\memory[11][4] ),
    .B(_05785_),
    .Y(_01204_)
  );
  NAND _09345_ (
    .A(\memory[29][4] ),
    .B(_05692_),
    .Y(_01205_)
  );
  NAND _09346_ (
    .A(\memory[10][4] ),
    .B(_05661_),
    .Y(_01206_)
  );
  NAND _09347_ (
    .A(\memory[27][4] ),
    .B(_05847_),
    .Y(_01207_)
  );
  NAND _09348_ (
    .A(\memory[8][4] ),
    .B(_05899_),
    .Y(_01208_)
  );
  NAND _09349_ (
    .A(\memory[26][4] ),
    .B(_05981_),
    .Y(_01209_)
  );
  NAND _09350_ (
    .A(\memory[6][4] ),
    .B(_06374_),
    .Y(_01210_)
  );
  NAND _09351_ (
    .A(\memory[18][4] ),
    .B(_05930_),
    .Y(_01211_)
  );
  NAND _09352_ (
    .A(\memory[13][4] ),
    .B(_06064_),
    .Y(_01212_)
  );
  NAND _09353_ (
    .A(\memory[16][4] ),
    .B(_05558_),
    .Y(_01213_)
  );
  NAND _09354_ (
    .A(\memory[5][4] ),
    .B(_05475_),
    .Y(_01214_)
  );
  NAND _09355_ (
    .A(\memory[0][4] ),
    .B(_06043_),
    .Y(_01215_)
  );
  NAND _09356_ (
    .A(\memory[9][4] ),
    .B(_06312_),
    .Y(_01216_)
  );
  NAND _09357_ (
    .A(\memory[30][4] ),
    .B(_06188_),
    .Y(_01217_)
  );
  NAND _09358_ (
    .A(\memory[15][4] ),
    .B(_06209_),
    .Y(_01218_)
  );
  NAND _09359_ (
    .A(\memory[31][4] ),
    .B(_06116_),
    .Y(_01219_)
  );
  NAND _09360_ (
    .A(\memory[3][4] ),
    .B(_06147_),
    .Y(_01220_)
  );
  NAND _09361_ (
    .A(\memory[19][4] ),
    .B(_06167_),
    .Y(_01221_)
  );
  NAND _09362_ (
    .A(\memory[22][4] ),
    .B(_06395_),
    .Y(_01222_)
  );
  NAND _09363_ (
    .A(\memory[14][4] ),
    .B(_06085_),
    .Y(_01223_)
  );
  NAND _09364_ (
    .A(\memory[23][4] ),
    .B(_06250_),
    .Y(_01224_)
  );
  NAND _09365_ (
    .A(\memory[2][4] ),
    .B(_05961_),
    .Y(_01225_)
  );
  NAND _09366_ (
    .A(\memory[7][4] ),
    .B(_06353_),
    .Y(_01226_)
  );
  NAND _09367_ (
    .A(\memory[24][4] ),
    .B(_06333_),
    .Y(_01227_)
  );
  NAND _09368_ (
    .A(\memory[25][4] ),
    .B(_06291_),
    .Y(_01228_)
  );
  AND _09369_ (
    .A(_01208_),
    .B(_01226_),
    .Y(_01229_)
  );
  AND _09370_ (
    .A(_01199_),
    .B(_01204_),
    .Y(_01230_)
  );
  AND _09371_ (
    .A(_01222_),
    .B(_01225_),
    .Y(_01231_)
  );
  AND _09372_ (
    .A(_01202_),
    .B(_01231_),
    .Y(_01232_)
  );
  AND _09373_ (
    .A(_01203_),
    .B(_01220_),
    .Y(_01233_)
  );
  AND _09374_ (
    .A(_01216_),
    .B(_01233_),
    .Y(_01234_)
  );
  AND _09375_ (
    .A(_01200_),
    .B(_01221_),
    .Y(_01235_)
  );
  AND _09376_ (
    .A(_01206_),
    .B(_01235_),
    .Y(_01236_)
  );
  AND _09377_ (
    .A(_01234_),
    .B(_01236_),
    .Y(_01237_)
  );
  AND _09378_ (
    .A(_01210_),
    .B(_01237_),
    .Y(_01238_)
  );
  AND _09379_ (
    .A(_01232_),
    .B(_01238_),
    .Y(_01239_)
  );
  AND _09380_ (
    .A(_01198_),
    .B(_01211_),
    .Y(_01240_)
  );
  AND _09381_ (
    .A(_01207_),
    .B(_01219_),
    .Y(_01241_)
  );
  AND _09382_ (
    .A(_01212_),
    .B(_01241_),
    .Y(_01242_)
  );
  AND _09383_ (
    .A(_01240_),
    .B(_01242_),
    .Y(_01243_)
  );
  AND _09384_ (
    .A(_01201_),
    .B(_01223_),
    .Y(_01244_)
  );
  AND _09385_ (
    .A(_01217_),
    .B(_01244_),
    .Y(_01245_)
  );
  AND _09386_ (
    .A(_01243_),
    .B(_01245_),
    .Y(_01246_)
  );
  AND _09387_ (
    .A(_01227_),
    .B(_01230_),
    .Y(_01247_)
  );
  AND _09388_ (
    .A(_01224_),
    .B(_01247_),
    .Y(_01248_)
  );
  AND _09389_ (
    .A(_01197_),
    .B(_01248_),
    .Y(_01249_)
  );
  AND _09390_ (
    .A(_01246_),
    .B(_01249_),
    .Y(_01250_)
  );
  AND _09391_ (
    .A(_01205_),
    .B(_01218_),
    .Y(_01251_)
  );
  AND _09392_ (
    .A(_01209_),
    .B(_01251_),
    .Y(_01252_)
  );
  AND _09393_ (
    .A(_01214_),
    .B(_01252_),
    .Y(_01253_)
  );
  AND _09394_ (
    .A(_01229_),
    .B(_01253_),
    .Y(_01254_)
  );
  AND _09395_ (
    .A(_01215_),
    .B(_01228_),
    .Y(_01255_)
  );
  AND _09396_ (
    .A(_01213_),
    .B(_01255_),
    .Y(_01256_)
  );
  AND _09397_ (
    .A(_01254_),
    .B(_01256_),
    .Y(_01257_)
  );
  AND _09398_ (
    .A(_01250_),
    .B(_01257_),
    .Y(_01258_)
  );
  NAND _09399_ (
    .A(_01239_),
    .B(_01258_),
    .Y(\data_mem_o[4] )
  );
  NAND _09400_ (
    .A(\memory[13][5] ),
    .B(_06064_),
    .Y(_01259_)
  );
  NAND _09401_ (
    .A(\memory[4][5] ),
    .B(_05733_),
    .Y(_01260_)
  );
  NAND _09402_ (
    .A(\memory[20][5] ),
    .B(_05806_),
    .Y(_01261_)
  );
  NAND _09403_ (
    .A(\memory[1][5] ),
    .B(_05599_),
    .Y(_01262_)
  );
  NAND _09404_ (
    .A(\memory[11][5] ),
    .B(_05785_),
    .Y(_01263_)
  );
  NAND _09405_ (
    .A(\memory[27][5] ),
    .B(_05847_),
    .Y(_01264_)
  );
  NAND _09406_ (
    .A(\memory[17][5] ),
    .B(_05754_),
    .Y(_01265_)
  );
  NAND _09407_ (
    .A(\memory[28][5] ),
    .B(_05826_),
    .Y(_01266_)
  );
  NAND _09408_ (
    .A(\memory[21][5] ),
    .B(_06023_),
    .Y(_01267_)
  );
  NAND _09409_ (
    .A(\memory[10][5] ),
    .B(_05661_),
    .Y(_01268_)
  );
  NAND _09410_ (
    .A(\memory[29][5] ),
    .B(_05692_),
    .Y(_01269_)
  );
  NAND _09411_ (
    .A(\memory[6][5] ),
    .B(_06374_),
    .Y(_01270_)
  );
  NAND _09412_ (
    .A(\memory[8][5] ),
    .B(_05899_),
    .Y(_01271_)
  );
  NAND _09413_ (
    .A(\memory[9][5] ),
    .B(_06312_),
    .Y(_01272_)
  );
  NAND _09414_ (
    .A(\memory[14][5] ),
    .B(_06085_),
    .Y(_01273_)
  );
  NAND _09415_ (
    .A(\memory[12][5] ),
    .B(_06002_),
    .Y(_01274_)
  );
  NAND _09416_ (
    .A(\memory[16][5] ),
    .B(_05558_),
    .Y(_01275_)
  );
  NAND _09417_ (
    .A(\memory[5][5] ),
    .B(_05475_),
    .Y(_01276_)
  );
  NAND _09418_ (
    .A(\memory[0][5] ),
    .B(_06043_),
    .Y(_01277_)
  );
  NAND _09419_ (
    .A(\memory[26][5] ),
    .B(_05981_),
    .Y(_01278_)
  );
  NAND _09420_ (
    .A(\memory[30][5] ),
    .B(_06188_),
    .Y(_01279_)
  );
  NAND _09421_ (
    .A(\memory[15][5] ),
    .B(_06209_),
    .Y(_01280_)
  );
  NAND _09422_ (
    .A(\memory[31][5] ),
    .B(_06116_),
    .Y(_01281_)
  );
  NAND _09423_ (
    .A(\memory[3][5] ),
    .B(_06147_),
    .Y(_01282_)
  );
  NAND _09424_ (
    .A(\memory[19][5] ),
    .B(_06167_),
    .Y(_01283_)
  );
  NAND _09425_ (
    .A(\memory[22][5] ),
    .B(_06395_),
    .Y(_01284_)
  );
  NAND _09426_ (
    .A(\memory[18][5] ),
    .B(_05930_),
    .Y(_01285_)
  );
  NAND _09427_ (
    .A(\memory[25][5] ),
    .B(_06291_),
    .Y(_01286_)
  );
  NAND _09428_ (
    .A(\memory[23][5] ),
    .B(_06250_),
    .Y(_01287_)
  );
  NAND _09429_ (
    .A(\memory[24][5] ),
    .B(_06333_),
    .Y(_01288_)
  );
  NAND _09430_ (
    .A(\memory[2][5] ),
    .B(_05961_),
    .Y(_01289_)
  );
  NAND _09431_ (
    .A(\memory[7][5] ),
    .B(_06353_),
    .Y(_01290_)
  );
  AND _09432_ (
    .A(_01263_),
    .B(_01274_),
    .Y(_01291_)
  );
  AND _09433_ (
    .A(_01271_),
    .B(_01290_),
    .Y(_01292_)
  );
  AND _09434_ (
    .A(_01265_),
    .B(_01285_),
    .Y(_01293_)
  );
  AND _09435_ (
    .A(_01284_),
    .B(_01289_),
    .Y(_01294_)
  );
  AND _09436_ (
    .A(_01262_),
    .B(_01294_),
    .Y(_01295_)
  );
  AND _09437_ (
    .A(_01260_),
    .B(_01282_),
    .Y(_01296_)
  );
  AND _09438_ (
    .A(_01272_),
    .B(_01296_),
    .Y(_01297_)
  );
  AND _09439_ (
    .A(_01261_),
    .B(_01283_),
    .Y(_01298_)
  );
  AND _09440_ (
    .A(_01268_),
    .B(_01298_),
    .Y(_01299_)
  );
  AND _09441_ (
    .A(_01297_),
    .B(_01299_),
    .Y(_01300_)
  );
  AND _09442_ (
    .A(_01270_),
    .B(_01300_),
    .Y(_01301_)
  );
  AND _09443_ (
    .A(_01295_),
    .B(_01301_),
    .Y(_01302_)
  );
  AND _09444_ (
    .A(_01264_),
    .B(_01281_),
    .Y(_01303_)
  );
  AND _09445_ (
    .A(_01259_),
    .B(_01303_),
    .Y(_01304_)
  );
  AND _09446_ (
    .A(_01266_),
    .B(_01273_),
    .Y(_01305_)
  );
  AND _09447_ (
    .A(_01279_),
    .B(_01305_),
    .Y(_01306_)
  );
  AND _09448_ (
    .A(_01304_),
    .B(_01306_),
    .Y(_01307_)
  );
  AND _09449_ (
    .A(_01267_),
    .B(_01287_),
    .Y(_01308_)
  );
  AND _09450_ (
    .A(_01288_),
    .B(_01291_),
    .Y(_01309_)
  );
  AND _09451_ (
    .A(_01308_),
    .B(_01309_),
    .Y(_01310_)
  );
  AND _09452_ (
    .A(_01293_),
    .B(_01310_),
    .Y(_01311_)
  );
  AND _09453_ (
    .A(_01307_),
    .B(_01311_),
    .Y(_01312_)
  );
  AND _09454_ (
    .A(_01269_),
    .B(_01280_),
    .Y(_01313_)
  );
  AND _09455_ (
    .A(_01278_),
    .B(_01313_),
    .Y(_01314_)
  );
  AND _09456_ (
    .A(_01276_),
    .B(_01314_),
    .Y(_01315_)
  );
  AND _09457_ (
    .A(_01292_),
    .B(_01315_),
    .Y(_01316_)
  );
  AND _09458_ (
    .A(_01277_),
    .B(_01286_),
    .Y(_01317_)
  );
  AND _09459_ (
    .A(_01275_),
    .B(_01317_),
    .Y(_01318_)
  );
  AND _09460_ (
    .A(_01316_),
    .B(_01318_),
    .Y(_01319_)
  );
  AND _09461_ (
    .A(_01312_),
    .B(_01319_),
    .Y(_01320_)
  );
  NAND _09462_ (
    .A(_01302_),
    .B(_01320_),
    .Y(\data_mem_o[5] )
  );
  NAND _09463_ (
    .A(\memory[13][6] ),
    .B(_06064_),
    .Y(_01321_)
  );
  NAND _09464_ (
    .A(\memory[4][6] ),
    .B(_05733_),
    .Y(_01322_)
  );
  NAND _09465_ (
    .A(\memory[20][6] ),
    .B(_05806_),
    .Y(_01323_)
  );
  NAND _09466_ (
    .A(\memory[1][6] ),
    .B(_05599_),
    .Y(_01324_)
  );
  NAND _09467_ (
    .A(\memory[11][6] ),
    .B(_05785_),
    .Y(_01325_)
  );
  NAND _09468_ (
    .A(\memory[27][6] ),
    .B(_05847_),
    .Y(_01326_)
  );
  NAND _09469_ (
    .A(\memory[17][6] ),
    .B(_05754_),
    .Y(_01327_)
  );
  NAND _09470_ (
    .A(\memory[28][6] ),
    .B(_05826_),
    .Y(_01328_)
  );
  NAND _09471_ (
    .A(\memory[21][6] ),
    .B(_06023_),
    .Y(_01329_)
  );
  NAND _09472_ (
    .A(\memory[10][6] ),
    .B(_05661_),
    .Y(_01330_)
  );
  NAND _09473_ (
    .A(\memory[29][6] ),
    .B(_05692_),
    .Y(_01331_)
  );
  NAND _09474_ (
    .A(\memory[6][6] ),
    .B(_06374_),
    .Y(_01332_)
  );
  NAND _09475_ (
    .A(\memory[8][6] ),
    .B(_05899_),
    .Y(_01333_)
  );
  NAND _09476_ (
    .A(\memory[9][6] ),
    .B(_06312_),
    .Y(_01334_)
  );
  NAND _09477_ (
    .A(\memory[14][6] ),
    .B(_06085_),
    .Y(_01335_)
  );
  NAND _09478_ (
    .A(\memory[12][6] ),
    .B(_06002_),
    .Y(_01336_)
  );
  NAND _09479_ (
    .A(\memory[16][6] ),
    .B(_05558_),
    .Y(_01337_)
  );
  NAND _09480_ (
    .A(\memory[5][6] ),
    .B(_05475_),
    .Y(_01338_)
  );
  NAND _09481_ (
    .A(\memory[0][6] ),
    .B(_06043_),
    .Y(_01339_)
  );
  NAND _09482_ (
    .A(\memory[26][6] ),
    .B(_05981_),
    .Y(_01340_)
  );
  NAND _09483_ (
    .A(\memory[30][6] ),
    .B(_06188_),
    .Y(_01341_)
  );
  NAND _09484_ (
    .A(\memory[15][6] ),
    .B(_06209_),
    .Y(_01342_)
  );
  NAND _09485_ (
    .A(\memory[31][6] ),
    .B(_06116_),
    .Y(_01343_)
  );
  NAND _09486_ (
    .A(\memory[3][6] ),
    .B(_06147_),
    .Y(_01344_)
  );
  NAND _09487_ (
    .A(\memory[19][6] ),
    .B(_06167_),
    .Y(_01345_)
  );
  NAND _09488_ (
    .A(\memory[22][6] ),
    .B(_06395_),
    .Y(_01346_)
  );
  NAND _09489_ (
    .A(\memory[18][6] ),
    .B(_05930_),
    .Y(_01347_)
  );
  NAND _09490_ (
    .A(\memory[25][6] ),
    .B(_06291_),
    .Y(_01348_)
  );
  NAND _09491_ (
    .A(\memory[23][6] ),
    .B(_06250_),
    .Y(_01349_)
  );
  NAND _09492_ (
    .A(\memory[24][6] ),
    .B(_06333_),
    .Y(_01350_)
  );
  NAND _09493_ (
    .A(\memory[2][6] ),
    .B(_05961_),
    .Y(_01351_)
  );
  NAND _09494_ (
    .A(\memory[7][6] ),
    .B(_06353_),
    .Y(_01352_)
  );
  AND _09495_ (
    .A(_01325_),
    .B(_01336_),
    .Y(_01353_)
  );
  AND _09496_ (
    .A(_01333_),
    .B(_01352_),
    .Y(_01354_)
  );
  AND _09497_ (
    .A(_01327_),
    .B(_01347_),
    .Y(_01355_)
  );
  AND _09498_ (
    .A(_01346_),
    .B(_01351_),
    .Y(_01356_)
  );
  AND _09499_ (
    .A(_01324_),
    .B(_01356_),
    .Y(_01357_)
  );
  AND _09500_ (
    .A(_01322_),
    .B(_01344_),
    .Y(_01358_)
  );
  AND _09501_ (
    .A(_01334_),
    .B(_01358_),
    .Y(_01359_)
  );
  AND _09502_ (
    .A(_01323_),
    .B(_01345_),
    .Y(_01360_)
  );
  AND _09503_ (
    .A(_01330_),
    .B(_01360_),
    .Y(_01361_)
  );
  AND _09504_ (
    .A(_01359_),
    .B(_01361_),
    .Y(_01362_)
  );
  AND _09505_ (
    .A(_01332_),
    .B(_01362_),
    .Y(_01363_)
  );
  AND _09506_ (
    .A(_01357_),
    .B(_01363_),
    .Y(_01364_)
  );
  AND _09507_ (
    .A(_01326_),
    .B(_01343_),
    .Y(_01365_)
  );
  AND _09508_ (
    .A(_01321_),
    .B(_01365_),
    .Y(_01366_)
  );
  AND _09509_ (
    .A(_01328_),
    .B(_01335_),
    .Y(_01367_)
  );
  AND _09510_ (
    .A(_01341_),
    .B(_01367_),
    .Y(_01368_)
  );
  AND _09511_ (
    .A(_01366_),
    .B(_01368_),
    .Y(_01369_)
  );
  AND _09512_ (
    .A(_01329_),
    .B(_01349_),
    .Y(_01370_)
  );
  AND _09513_ (
    .A(_01350_),
    .B(_01353_),
    .Y(_01371_)
  );
  AND _09514_ (
    .A(_01370_),
    .B(_01371_),
    .Y(_01372_)
  );
  AND _09515_ (
    .A(_01355_),
    .B(_01372_),
    .Y(_01373_)
  );
  AND _09516_ (
    .A(_01369_),
    .B(_01373_),
    .Y(_01374_)
  );
  AND _09517_ (
    .A(_01331_),
    .B(_01342_),
    .Y(_01375_)
  );
  AND _09518_ (
    .A(_01340_),
    .B(_01375_),
    .Y(_01376_)
  );
  AND _09519_ (
    .A(_01338_),
    .B(_01376_),
    .Y(_01377_)
  );
  AND _09520_ (
    .A(_01354_),
    .B(_01377_),
    .Y(_01378_)
  );
  AND _09521_ (
    .A(_01339_),
    .B(_01348_),
    .Y(_01379_)
  );
  AND _09522_ (
    .A(_01337_),
    .B(_01379_),
    .Y(_01380_)
  );
  AND _09523_ (
    .A(_01378_),
    .B(_01380_),
    .Y(_01381_)
  );
  AND _09524_ (
    .A(_01374_),
    .B(_01381_),
    .Y(_01382_)
  );
  NAND _09525_ (
    .A(_01364_),
    .B(_01382_),
    .Y(\data_mem_o[6] )
  );
  NAND _09526_ (
    .A(\memory[0][7] ),
    .B(_06043_),
    .Y(_01383_)
  );
  NAND _09527_ (
    .A(\memory[4][7] ),
    .B(_05733_),
    .Y(_01384_)
  );
  NAND _09528_ (
    .A(\memory[17][7] ),
    .B(_05754_),
    .Y(_01385_)
  );
  NAND _09529_ (
    .A(\memory[1][7] ),
    .B(_05599_),
    .Y(_01386_)
  );
  NAND _09530_ (
    .A(\memory[20][7] ),
    .B(_05806_),
    .Y(_01387_)
  );
  NAND _09531_ (
    .A(\memory[5][7] ),
    .B(_05475_),
    .Y(_01388_)
  );
  NAND _09532_ (
    .A(\memory[29][7] ),
    .B(_05692_),
    .Y(_01389_)
  );
  NAND _09533_ (
    .A(\memory[16][7] ),
    .B(_05558_),
    .Y(_01390_)
  );
  NAND _09534_ (
    .A(\memory[28][7] ),
    .B(_05826_),
    .Y(_01391_)
  );
  NAND _09535_ (
    .A(\memory[10][7] ),
    .B(_05661_),
    .Y(_01392_)
  );
  NAND _09536_ (
    .A(\memory[27][7] ),
    .B(_05847_),
    .Y(_01393_)
  );
  NAND _09537_ (
    .A(\memory[22][7] ),
    .B(_06395_),
    .Y(_01394_)
  );
  NAND _09538_ (
    .A(\memory[2][7] ),
    .B(_05961_),
    .Y(_01395_)
  );
  AND _09539_ (
    .A(_01394_),
    .B(_01395_),
    .Y(_01396_)
  );
  NAND _09540_ (
    .A(\memory[7][7] ),
    .B(_06353_),
    .Y(_01397_)
  );
  NAND _09541_ (
    .A(\memory[23][7] ),
    .B(_06250_),
    .Y(_01398_)
  );
  NAND _09542_ (
    .A(\memory[13][7] ),
    .B(_06064_),
    .Y(_01399_)
  );
  NAND _09543_ (
    .A(\memory[12][7] ),
    .B(_06002_),
    .Y(_01400_)
  );
  NAND _09544_ (
    .A(\memory[21][7] ),
    .B(_06023_),
    .Y(_01401_)
  );
  NAND _09545_ (
    .A(\memory[11][7] ),
    .B(_05785_),
    .Y(_01402_)
  );
  NAND _09546_ (
    .A(\memory[25][7] ),
    .B(_06291_),
    .Y(_01403_)
  );
  NAND _09547_ (
    .A(\memory[31][7] ),
    .B(_06116_),
    .Y(_01404_)
  );
  NAND _09548_ (
    .A(\memory[3][7] ),
    .B(_06147_),
    .Y(_01405_)
  );
  NAND _09549_ (
    .A(\memory[19][7] ),
    .B(_06167_),
    .Y(_01406_)
  );
  NAND _09550_ (
    .A(\memory[15][7] ),
    .B(_06209_),
    .Y(_01407_)
  );
  NAND _09551_ (
    .A(\memory[30][7] ),
    .B(_06188_),
    .Y(_01408_)
  );
  NAND _09552_ (
    .A(\memory[8][7] ),
    .B(_05899_),
    .Y(_01409_)
  );
  NAND _09553_ (
    .A(\memory[6][7] ),
    .B(_06374_),
    .Y(_01410_)
  );
  NAND _09554_ (
    .A(\memory[9][7] ),
    .B(_06312_),
    .Y(_01411_)
  );
  NAND _09555_ (
    .A(\memory[26][7] ),
    .B(_05981_),
    .Y(_01412_)
  );
  NAND _09556_ (
    .A(\memory[14][7] ),
    .B(_06085_),
    .Y(_01413_)
  );
  NAND _09557_ (
    .A(\memory[18][7] ),
    .B(_05930_),
    .Y(_01414_)
  );
  NAND _09558_ (
    .A(\memory[24][7] ),
    .B(_06333_),
    .Y(_01415_)
  );
  AND _09559_ (
    .A(_01400_),
    .B(_01402_),
    .Y(_01416_)
  );
  AND _09560_ (
    .A(_01397_),
    .B(_01409_),
    .Y(_01417_)
  );
  AND _09561_ (
    .A(_01389_),
    .B(_01407_),
    .Y(_01418_)
  );
  AND _09562_ (
    .A(_01412_),
    .B(_01418_),
    .Y(_01419_)
  );
  AND _09563_ (
    .A(_01388_),
    .B(_01419_),
    .Y(_01420_)
  );
  AND _09564_ (
    .A(_01417_),
    .B(_01420_),
    .Y(_01421_)
  );
  AND _09565_ (
    .A(_01383_),
    .B(_01403_),
    .Y(_01422_)
  );
  AND _09566_ (
    .A(_01390_),
    .B(_01422_),
    .Y(_01423_)
  );
  AND _09567_ (
    .A(_01421_),
    .B(_01423_),
    .Y(_01424_)
  );
  AND _09568_ (
    .A(_01386_),
    .B(_01396_),
    .Y(_01425_)
  );
  AND _09569_ (
    .A(_01384_),
    .B(_01405_),
    .Y(_01426_)
  );
  AND _09570_ (
    .A(_01411_),
    .B(_01426_),
    .Y(_01427_)
  );
  AND _09571_ (
    .A(_01387_),
    .B(_01406_),
    .Y(_01428_)
  );
  AND _09572_ (
    .A(_01392_),
    .B(_01428_),
    .Y(_01429_)
  );
  AND _09573_ (
    .A(_01427_),
    .B(_01429_),
    .Y(_01430_)
  );
  AND _09574_ (
    .A(_01410_),
    .B(_01430_),
    .Y(_01431_)
  );
  AND _09575_ (
    .A(_01425_),
    .B(_01431_),
    .Y(_01432_)
  );
  AND _09576_ (
    .A(_01424_),
    .B(_01432_),
    .Y(_01433_)
  );
  AND _09577_ (
    .A(_01385_),
    .B(_01414_),
    .Y(_01434_)
  );
  AND _09578_ (
    .A(_01393_),
    .B(_01404_),
    .Y(_01435_)
  );
  AND _09579_ (
    .A(_01399_),
    .B(_01435_),
    .Y(_01436_)
  );
  AND _09580_ (
    .A(_01434_),
    .B(_01436_),
    .Y(_01437_)
  );
  AND _09581_ (
    .A(_01391_),
    .B(_01413_),
    .Y(_01438_)
  );
  AND _09582_ (
    .A(_01408_),
    .B(_01438_),
    .Y(_01439_)
  );
  AND _09583_ (
    .A(_01415_),
    .B(_01416_),
    .Y(_01440_)
  );
  AND _09584_ (
    .A(_01398_),
    .B(_01440_),
    .Y(_01441_)
  );
  AND _09585_ (
    .A(_01401_),
    .B(_01441_),
    .Y(_01442_)
  );
  AND _09586_ (
    .A(_01439_),
    .B(_01442_),
    .Y(_01443_)
  );
  AND _09587_ (
    .A(_01437_),
    .B(_01443_),
    .Y(_01444_)
  );
  NAND _09588_ (
    .A(_01433_),
    .B(_01444_),
    .Y(\data_mem_o[7] )
  );
  NOR _09589_ (
    .A(\addr_i[3] ),
    .B(\addr_i[2] ),
    .Y(_01445_)
  );
  NOR _09590_ (
    .A(\addr_i[1] ),
    .B(\addr_i[0] ),
    .Y(_01446_)
  );
  AND _09591_ (
    .A(_05351_),
    .B(_01446_),
    .Y(_01447_)
  );
  AND _09592_ (
    .A(_05351_),
    .B(_01445_),
    .Y(_01448_)
  );
  AND _09593_ (
    .A(_01445_),
    .B(_01447_),
    .Y(_01449_)
  );
  NAND _09594_ (
    .A(_01445_),
    .B(_01447_),
    .Y(_01450_)
  );
  NAND _09595_ (
    .A(\memory[0][0] ),
    .B(_01449_),
    .Y(_01451_)
  );
  AND _09596_ (
    .A(\addr_i[1] ),
    .B(_05330_),
    .Y(_01452_)
  );
  AND _09597_ (
    .A(_01448_),
    .B(_01452_),
    .Y(_01453_)
  );
  NAND _09598_ (
    .A(_01448_),
    .B(_01452_),
    .Y(_01454_)
  );
  NAND _09599_ (
    .A(\memory[2][0] ),
    .B(_01453_),
    .Y(_01455_)
  );
  AND _09600_ (
    .A(_01451_),
    .B(_01455_),
    .Y(_01456_)
  );
  AND _09601_ (
    .A(\addr_i[3] ),
    .B(\addr_i[2] ),
    .Y(_01457_)
  );
  AND _09602_ (
    .A(_01447_),
    .B(_01457_),
    .Y(_01458_)
  );
  NAND _09603_ (
    .A(_01447_),
    .B(_01457_),
    .Y(_01459_)
  );
  NAND _09604_ (
    .A(\memory[12][0] ),
    .B(_01458_),
    .Y(_01460_)
  );
  AND _09605_ (
    .A(\addr_i[4] ),
    .B(_01446_),
    .Y(_01461_)
  );
  AND _09606_ (
    .A(_01457_),
    .B(_01461_),
    .Y(_01462_)
  );
  NAND _09607_ (
    .A(_01457_),
    .B(_01461_),
    .Y(_01463_)
  );
  NAND _09608_ (
    .A(\memory[28][0] ),
    .B(_01462_),
    .Y(_01464_)
  );
  AND _09609_ (
    .A(_01460_),
    .B(_01464_),
    .Y(_01465_)
  );
  AND _09610_ (
    .A(_01456_),
    .B(_01465_),
    .Y(_01466_)
  );
  AND _09611_ (
    .A(_05341_),
    .B(\addr_i[2] ),
    .Y(_01467_)
  );
  AND _09612_ (
    .A(_01452_),
    .B(_01467_),
    .Y(_01468_)
  );
  AND _09613_ (
    .A(\addr_i[4] ),
    .B(_01468_),
    .Y(_01469_)
  );
  NAND _09614_ (
    .A(\addr_i[4] ),
    .B(_01468_),
    .Y(_01470_)
  );
  NAND _09615_ (
    .A(\memory[22][0] ),
    .B(_01469_),
    .Y(_01471_)
  );
  NOR _09616_ (
    .A(\addr_i[1] ),
    .B(_05330_),
    .Y(_01472_)
  );
  AND _09617_ (
    .A(_01467_),
    .B(_01472_),
    .Y(_01473_)
  );
  AND _09618_ (
    .A(\addr_i[4] ),
    .B(_01473_),
    .Y(_01474_)
  );
  NAND _09619_ (
    .A(\addr_i[4] ),
    .B(_01473_),
    .Y(_01475_)
  );
  NAND _09620_ (
    .A(\memory[21][0] ),
    .B(_01474_),
    .Y(_01476_)
  );
  AND _09621_ (
    .A(_01471_),
    .B(_01476_),
    .Y(_01477_)
  );
  AND _09622_ (
    .A(\addr_i[4] ),
    .B(_01445_),
    .Y(_01478_)
  );
  AND _09623_ (
    .A(_01472_),
    .B(_01478_),
    .Y(_01479_)
  );
  NAND _09624_ (
    .A(_01472_),
    .B(_01478_),
    .Y(_01480_)
  );
  NAND _09625_ (
    .A(\memory[17][0] ),
    .B(_01479_),
    .Y(_01481_)
  );
  NOR _09626_ (
    .A(_05341_),
    .B(\addr_i[2] ),
    .Y(_01482_)
  );
  AND _09627_ (
    .A(_01452_),
    .B(_01482_),
    .Y(_01483_)
  );
  AND _09628_ (
    .A(\addr_i[4] ),
    .B(_01483_),
    .Y(_01484_)
  );
  NAND _09629_ (
    .A(\addr_i[4] ),
    .B(_01483_),
    .Y(_01485_)
  );
  NAND _09630_ (
    .A(\memory[26][0] ),
    .B(_01484_),
    .Y(_01486_)
  );
  AND _09631_ (
    .A(_01481_),
    .B(_01486_),
    .Y(_01487_)
  );
  AND _09632_ (
    .A(_01477_),
    .B(_01487_),
    .Y(_01488_)
  );
  AND _09633_ (
    .A(_01466_),
    .B(_01488_),
    .Y(_01489_)
  );
  AND _09634_ (
    .A(_01452_),
    .B(_01457_),
    .Y(_01490_)
  );
  AND _09635_ (
    .A(\addr_i[4] ),
    .B(_01490_),
    .Y(_01491_)
  );
  NAND _09636_ (
    .A(\addr_i[4] ),
    .B(_01490_),
    .Y(_01492_)
  );
  NAND _09637_ (
    .A(\memory[30][0] ),
    .B(_01491_),
    .Y(_01493_)
  );
  AND _09638_ (
    .A(_01472_),
    .B(_01482_),
    .Y(_01494_)
  );
  AND _09639_ (
    .A(_05351_),
    .B(_01494_),
    .Y(_01495_)
  );
  NAND _09640_ (
    .A(_05351_),
    .B(_01494_),
    .Y(_01496_)
  );
  NAND _09641_ (
    .A(\memory[9][0] ),
    .B(_01495_),
    .Y(_01497_)
  );
  AND _09642_ (
    .A(_01493_),
    .B(_01497_),
    .Y(_01498_)
  );
  AND _09643_ (
    .A(\addr_i[1] ),
    .B(\addr_i[0] ),
    .Y(_01499_)
  );
  AND _09644_ (
    .A(_01457_),
    .B(_01499_),
    .Y(_01500_)
  );
  AND _09645_ (
    .A(_05351_),
    .B(_01500_),
    .Y(_01501_)
  );
  NAND _09646_ (
    .A(_05351_),
    .B(_01500_),
    .Y(_01502_)
  );
  NAND _09647_ (
    .A(\memory[15][0] ),
    .B(_01501_),
    .Y(_01503_)
  );
  AND _09648_ (
    .A(\addr_i[4] ),
    .B(_01500_),
    .Y(_01504_)
  );
  NAND _09649_ (
    .A(\addr_i[4] ),
    .B(_01500_),
    .Y(_01505_)
  );
  NAND _09650_ (
    .A(\memory[31][0] ),
    .B(_01504_),
    .Y(_01506_)
  );
  AND _09651_ (
    .A(_01503_),
    .B(_01506_),
    .Y(_01507_)
  );
  AND _09652_ (
    .A(_01498_),
    .B(_01507_),
    .Y(_01508_)
  );
  AND _09653_ (
    .A(_01457_),
    .B(_01472_),
    .Y(_01509_)
  );
  AND _09654_ (
    .A(\addr_i[4] ),
    .B(_01509_),
    .Y(_01510_)
  );
  NAND _09655_ (
    .A(\addr_i[4] ),
    .B(_01509_),
    .Y(_01511_)
  );
  NAND _09656_ (
    .A(\memory[29][0] ),
    .B(_01510_),
    .Y(_01512_)
  );
  AND _09657_ (
    .A(_01448_),
    .B(_01499_),
    .Y(_01513_)
  );
  NAND _09658_ (
    .A(_01448_),
    .B(_01499_),
    .Y(_01514_)
  );
  NAND _09659_ (
    .A(\memory[3][0] ),
    .B(_01513_),
    .Y(_01515_)
  );
  AND _09660_ (
    .A(_01512_),
    .B(_01515_),
    .Y(_01516_)
  );
  AND _09661_ (
    .A(_05351_),
    .B(_01468_),
    .Y(_01517_)
  );
  NAND _09662_ (
    .A(_05351_),
    .B(_01468_),
    .Y(_01518_)
  );
  NAND _09663_ (
    .A(\memory[6][0] ),
    .B(_01517_),
    .Y(_01519_)
  );
  AND _09664_ (
    .A(_05351_),
    .B(_01509_),
    .Y(_01520_)
  );
  NAND _09665_ (
    .A(_05351_),
    .B(_01509_),
    .Y(_01521_)
  );
  NAND _09666_ (
    .A(\memory[13][0] ),
    .B(_01520_),
    .Y(_01522_)
  );
  AND _09667_ (
    .A(_01519_),
    .B(_01522_),
    .Y(_01523_)
  );
  AND _09668_ (
    .A(_01516_),
    .B(_01523_),
    .Y(_01524_)
  );
  AND _09669_ (
    .A(_01508_),
    .B(_01524_),
    .Y(_01525_)
  );
  AND _09670_ (
    .A(_01489_),
    .B(_01525_),
    .Y(_01526_)
  );
  AND _09671_ (
    .A(_01447_),
    .B(_01482_),
    .Y(_01527_)
  );
  NAND _09672_ (
    .A(_01447_),
    .B(_01482_),
    .Y(_01528_)
  );
  NAND _09673_ (
    .A(\memory[8][0] ),
    .B(_01527_),
    .Y(_01529_)
  );
  AND _09674_ (
    .A(_01447_),
    .B(_01467_),
    .Y(_01530_)
  );
  NAND _09675_ (
    .A(_01447_),
    .B(_01467_),
    .Y(_01531_)
  );
  NAND _09676_ (
    .A(\memory[4][0] ),
    .B(_01530_),
    .Y(_01532_)
  );
  AND _09677_ (
    .A(_01529_),
    .B(_01532_),
    .Y(_01533_)
  );
  AND _09678_ (
    .A(_01478_),
    .B(_01499_),
    .Y(_01534_)
  );
  NAND _09679_ (
    .A(_01478_),
    .B(_01499_),
    .Y(_01535_)
  );
  NAND _09680_ (
    .A(\memory[19][0] ),
    .B(_01534_),
    .Y(_01536_)
  );
  AND _09681_ (
    .A(_01467_),
    .B(_01499_),
    .Y(_01537_)
  );
  AND _09682_ (
    .A(_05351_),
    .B(_01537_),
    .Y(_01538_)
  );
  NAND _09683_ (
    .A(_05351_),
    .B(_01537_),
    .Y(_01539_)
  );
  NAND _09684_ (
    .A(\memory[7][0] ),
    .B(_01538_),
    .Y(_01540_)
  );
  AND _09685_ (
    .A(_01536_),
    .B(_01540_),
    .Y(_01541_)
  );
  AND _09686_ (
    .A(_01533_),
    .B(_01541_),
    .Y(_01542_)
  );
  AND _09687_ (
    .A(_05351_),
    .B(_01490_),
    .Y(_01543_)
  );
  NAND _09688_ (
    .A(_05351_),
    .B(_01490_),
    .Y(_01544_)
  );
  NAND _09689_ (
    .A(\memory[14][0] ),
    .B(_01543_),
    .Y(_01545_)
  );
  AND _09690_ (
    .A(\addr_i[4] ),
    .B(_01537_),
    .Y(_01546_)
  );
  NAND _09691_ (
    .A(\addr_i[4] ),
    .B(_01537_),
    .Y(_01547_)
  );
  NAND _09692_ (
    .A(\memory[23][0] ),
    .B(_01546_),
    .Y(_01548_)
  );
  AND _09693_ (
    .A(_01545_),
    .B(_01548_),
    .Y(_01549_)
  );
  AND _09694_ (
    .A(_01461_),
    .B(_01482_),
    .Y(_01550_)
  );
  NAND _09695_ (
    .A(_01461_),
    .B(_01482_),
    .Y(_01551_)
  );
  NAND _09696_ (
    .A(\memory[24][0] ),
    .B(_01550_),
    .Y(_01552_)
  );
  AND _09697_ (
    .A(_01461_),
    .B(_01467_),
    .Y(_01553_)
  );
  NAND _09698_ (
    .A(_01461_),
    .B(_01467_),
    .Y(_01554_)
  );
  NAND _09699_ (
    .A(\memory[20][0] ),
    .B(_01553_),
    .Y(_01555_)
  );
  AND _09700_ (
    .A(_01552_),
    .B(_01555_),
    .Y(_01556_)
  );
  AND _09701_ (
    .A(_01549_),
    .B(_01556_),
    .Y(_01557_)
  );
  AND _09702_ (
    .A(_01542_),
    .B(_01557_),
    .Y(_01558_)
  );
  AND _09703_ (
    .A(\addr_i[4] ),
    .B(_01494_),
    .Y(_01559_)
  );
  NAND _09704_ (
    .A(\addr_i[4] ),
    .B(_01494_),
    .Y(_01560_)
  );
  NAND _09705_ (
    .A(\memory[25][0] ),
    .B(_01559_),
    .Y(_01561_)
  );
  AND _09706_ (
    .A(_01482_),
    .B(_01499_),
    .Y(_01562_)
  );
  AND _09707_ (
    .A(\addr_i[4] ),
    .B(_01562_),
    .Y(_01563_)
  );
  NAND _09708_ (
    .A(\addr_i[4] ),
    .B(_01562_),
    .Y(_01564_)
  );
  NAND _09709_ (
    .A(\memory[27][0] ),
    .B(_01563_),
    .Y(_01565_)
  );
  AND _09710_ (
    .A(_01561_),
    .B(_01565_),
    .Y(_01566_)
  );
  AND _09711_ (
    .A(_01446_),
    .B(_01478_),
    .Y(_01567_)
  );
  NAND _09712_ (
    .A(_01446_),
    .B(_01478_),
    .Y(_01568_)
  );
  NAND _09713_ (
    .A(\memory[16][0] ),
    .B(_01567_),
    .Y(_01569_)
  );
  AND _09714_ (
    .A(_01448_),
    .B(_01472_),
    .Y(_01570_)
  );
  NAND _09715_ (
    .A(_01448_),
    .B(_01472_),
    .Y(_01571_)
  );
  NAND _09716_ (
    .A(\memory[1][0] ),
    .B(_01570_),
    .Y(_01572_)
  );
  AND _09717_ (
    .A(_01569_),
    .B(_01572_),
    .Y(_01573_)
  );
  AND _09718_ (
    .A(_01566_),
    .B(_01573_),
    .Y(_01574_)
  );
  AND _09719_ (
    .A(_05351_),
    .B(_01562_),
    .Y(_01575_)
  );
  NAND _09720_ (
    .A(_05351_),
    .B(_01562_),
    .Y(_01576_)
  );
  NAND _09721_ (
    .A(\memory[11][0] ),
    .B(_01575_),
    .Y(_01577_)
  );
  AND _09722_ (
    .A(_05351_),
    .B(_01483_),
    .Y(_01578_)
  );
  NAND _09723_ (
    .A(_05351_),
    .B(_01483_),
    .Y(_01579_)
  );
  NAND _09724_ (
    .A(\memory[10][0] ),
    .B(_01578_),
    .Y(_01580_)
  );
  AND _09725_ (
    .A(_01577_),
    .B(_01580_),
    .Y(_01581_)
  );
  AND _09726_ (
    .A(_01452_),
    .B(_01478_),
    .Y(_01582_)
  );
  NAND _09727_ (
    .A(_01452_),
    .B(_01478_),
    .Y(_01583_)
  );
  NAND _09728_ (
    .A(\memory[18][0] ),
    .B(_01582_),
    .Y(_01584_)
  );
  AND _09729_ (
    .A(_05351_),
    .B(_01473_),
    .Y(_01585_)
  );
  NAND _09730_ (
    .A(_05351_),
    .B(_01473_),
    .Y(_01586_)
  );
  NAND _09731_ (
    .A(\memory[5][0] ),
    .B(_01585_),
    .Y(_01587_)
  );
  AND _09732_ (
    .A(_01584_),
    .B(_01587_),
    .Y(_01588_)
  );
  AND _09733_ (
    .A(_01581_),
    .B(_01588_),
    .Y(_01589_)
  );
  AND _09734_ (
    .A(_01574_),
    .B(_01589_),
    .Y(_01590_)
  );
  AND _09735_ (
    .A(_01558_),
    .B(_01590_),
    .Y(_01591_)
  );
  NAND _09736_ (
    .A(_01526_),
    .B(_01591_),
    .Y(_01592_)
  );
  AND _09737_ (
    .A(MemRead_i),
    .B(_01592_),
    .Y(\data_o[0] )
  );
  NAND _09738_ (
    .A(\memory[22][1] ),
    .B(_01469_),
    .Y(_01593_)
  );
  NAND _09739_ (
    .A(\memory[4][1] ),
    .B(_01530_),
    .Y(_01594_)
  );
  AND _09740_ (
    .A(_01593_),
    .B(_01594_),
    .Y(_01595_)
  );
  NAND _09741_ (
    .A(\memory[6][1] ),
    .B(_01517_),
    .Y(_01596_)
  );
  NAND _09742_ (
    .A(\memory[7][1] ),
    .B(_01538_),
    .Y(_01597_)
  );
  AND _09743_ (
    .A(_01596_),
    .B(_01597_),
    .Y(_01598_)
  );
  AND _09744_ (
    .A(_01595_),
    .B(_01598_),
    .Y(_01599_)
  );
  NAND _09745_ (
    .A(\memory[8][1] ),
    .B(_01527_),
    .Y(_01600_)
  );
  NAND _09746_ (
    .A(\memory[27][1] ),
    .B(_01563_),
    .Y(_01601_)
  );
  AND _09747_ (
    .A(_01600_),
    .B(_01601_),
    .Y(_01602_)
  );
  NAND _09748_ (
    .A(\memory[31][1] ),
    .B(_01504_),
    .Y(_01603_)
  );
  NAND _09749_ (
    .A(\memory[25][1] ),
    .B(_01559_),
    .Y(_01604_)
  );
  AND _09750_ (
    .A(_01603_),
    .B(_01604_),
    .Y(_01605_)
  );
  AND _09751_ (
    .A(_01602_),
    .B(_01605_),
    .Y(_01606_)
  );
  AND _09752_ (
    .A(_01599_),
    .B(_01606_),
    .Y(_01607_)
  );
  NAND _09753_ (
    .A(\memory[12][1] ),
    .B(_01458_),
    .Y(_01608_)
  );
  NAND _09754_ (
    .A(\memory[30][1] ),
    .B(_01491_),
    .Y(_01609_)
  );
  AND _09755_ (
    .A(_01608_),
    .B(_01609_),
    .Y(_01610_)
  );
  NAND _09756_ (
    .A(\memory[13][1] ),
    .B(_01520_),
    .Y(_01611_)
  );
  NAND _09757_ (
    .A(\memory[26][1] ),
    .B(_01484_),
    .Y(_01612_)
  );
  AND _09758_ (
    .A(_01611_),
    .B(_01612_),
    .Y(_01613_)
  );
  AND _09759_ (
    .A(_01610_),
    .B(_01613_),
    .Y(_01614_)
  );
  NAND _09760_ (
    .A(\memory[20][1] ),
    .B(_01553_),
    .Y(_01615_)
  );
  NAND _09761_ (
    .A(\memory[11][1] ),
    .B(_01575_),
    .Y(_01616_)
  );
  AND _09762_ (
    .A(_01615_),
    .B(_01616_),
    .Y(_01617_)
  );
  NAND _09763_ (
    .A(\memory[0][1] ),
    .B(_01449_),
    .Y(_01618_)
  );
  NAND _09764_ (
    .A(\memory[9][1] ),
    .B(_01495_),
    .Y(_01619_)
  );
  AND _09765_ (
    .A(_01618_),
    .B(_01619_),
    .Y(_01620_)
  );
  AND _09766_ (
    .A(_01617_),
    .B(_01620_),
    .Y(_01621_)
  );
  AND _09767_ (
    .A(_01614_),
    .B(_01621_),
    .Y(_01622_)
  );
  AND _09768_ (
    .A(_01607_),
    .B(_01622_),
    .Y(_01623_)
  );
  NAND _09769_ (
    .A(\memory[10][1] ),
    .B(_01578_),
    .Y(_01624_)
  );
  NAND _09770_ (
    .A(\memory[16][1] ),
    .B(_01567_),
    .Y(_01625_)
  );
  AND _09771_ (
    .A(_01624_),
    .B(_01625_),
    .Y(_01626_)
  );
  NAND _09772_ (
    .A(\memory[1][1] ),
    .B(_01570_),
    .Y(_01627_)
  );
  NAND _09773_ (
    .A(\memory[15][1] ),
    .B(_01501_),
    .Y(_01628_)
  );
  AND _09774_ (
    .A(_01627_),
    .B(_01628_),
    .Y(_01629_)
  );
  AND _09775_ (
    .A(_01626_),
    .B(_01629_),
    .Y(_01630_)
  );
  NAND _09776_ (
    .A(\memory[17][1] ),
    .B(_01479_),
    .Y(_01631_)
  );
  NAND _09777_ (
    .A(\memory[18][1] ),
    .B(_01582_),
    .Y(_01632_)
  );
  AND _09778_ (
    .A(_01631_),
    .B(_01632_),
    .Y(_01633_)
  );
  NAND _09779_ (
    .A(\memory[19][1] ),
    .B(_01534_),
    .Y(_01634_)
  );
  NAND _09780_ (
    .A(\memory[28][1] ),
    .B(_01462_),
    .Y(_01635_)
  );
  AND _09781_ (
    .A(_01634_),
    .B(_01635_),
    .Y(_01636_)
  );
  AND _09782_ (
    .A(_01633_),
    .B(_01636_),
    .Y(_01637_)
  );
  AND _09783_ (
    .A(_01630_),
    .B(_01637_),
    .Y(_01638_)
  );
  NAND _09784_ (
    .A(\memory[23][1] ),
    .B(_01546_),
    .Y(_01639_)
  );
  NAND _09785_ (
    .A(\memory[24][1] ),
    .B(_01550_),
    .Y(_01640_)
  );
  AND _09786_ (
    .A(_01639_),
    .B(_01640_),
    .Y(_01641_)
  );
  NAND _09787_ (
    .A(\memory[2][1] ),
    .B(_01453_),
    .Y(_01642_)
  );
  NAND _09788_ (
    .A(\memory[3][1] ),
    .B(_01513_),
    .Y(_01643_)
  );
  AND _09789_ (
    .A(_01642_),
    .B(_01643_),
    .Y(_01644_)
  );
  AND _09790_ (
    .A(_01641_),
    .B(_01644_),
    .Y(_01645_)
  );
  NAND _09791_ (
    .A(\memory[14][1] ),
    .B(_01543_),
    .Y(_01646_)
  );
  NAND _09792_ (
    .A(\memory[21][1] ),
    .B(_01474_),
    .Y(_01647_)
  );
  AND _09793_ (
    .A(_01646_),
    .B(_01647_),
    .Y(_01648_)
  );
  NAND _09794_ (
    .A(\memory[29][1] ),
    .B(_01510_),
    .Y(_01649_)
  );
  NAND _09795_ (
    .A(\memory[5][1] ),
    .B(_01585_),
    .Y(_01650_)
  );
  AND _09796_ (
    .A(_01649_),
    .B(_01650_),
    .Y(_01651_)
  );
  AND _09797_ (
    .A(_01648_),
    .B(_01651_),
    .Y(_01652_)
  );
  AND _09798_ (
    .A(_01645_),
    .B(_01652_),
    .Y(_01653_)
  );
  AND _09799_ (
    .A(_01638_),
    .B(_01653_),
    .Y(_01654_)
  );
  NAND _09800_ (
    .A(_01623_),
    .B(_01654_),
    .Y(_01655_)
  );
  AND _09801_ (
    .A(MemRead_i),
    .B(_01655_),
    .Y(\data_o[1] )
  );
  NAND _09802_ (
    .A(\memory[29][2] ),
    .B(_01510_),
    .Y(_01656_)
  );
  NAND _09803_ (
    .A(\memory[0][2] ),
    .B(_01449_),
    .Y(_01657_)
  );
  AND _09804_ (
    .A(_01656_),
    .B(_01657_),
    .Y(_01658_)
  );
  NAND _09805_ (
    .A(\memory[19][2] ),
    .B(_01534_),
    .Y(_01659_)
  );
  NAND _09806_ (
    .A(\memory[28][2] ),
    .B(_01462_),
    .Y(_01660_)
  );
  AND _09807_ (
    .A(_01659_),
    .B(_01660_),
    .Y(_01661_)
  );
  AND _09808_ (
    .A(_01658_),
    .B(_01661_),
    .Y(_01662_)
  );
  NAND _09809_ (
    .A(\memory[7][2] ),
    .B(_01538_),
    .Y(_01663_)
  );
  NAND _09810_ (
    .A(\memory[4][2] ),
    .B(_01530_),
    .Y(_01664_)
  );
  AND _09811_ (
    .A(_01663_),
    .B(_01664_),
    .Y(_01665_)
  );
  NAND _09812_ (
    .A(\memory[11][2] ),
    .B(_01575_),
    .Y(_01666_)
  );
  NAND _09813_ (
    .A(\memory[9][2] ),
    .B(_01495_),
    .Y(_01667_)
  );
  AND _09814_ (
    .A(_01666_),
    .B(_01667_),
    .Y(_01668_)
  );
  AND _09815_ (
    .A(_01665_),
    .B(_01668_),
    .Y(_01669_)
  );
  AND _09816_ (
    .A(_01662_),
    .B(_01669_),
    .Y(_01670_)
  );
  NAND _09817_ (
    .A(\memory[15][2] ),
    .B(_01501_),
    .Y(_01671_)
  );
  NAND _09818_ (
    .A(\memory[26][2] ),
    .B(_01484_),
    .Y(_01672_)
  );
  AND _09819_ (
    .A(_01671_),
    .B(_01672_),
    .Y(_01673_)
  );
  NAND _09820_ (
    .A(\memory[2][2] ),
    .B(_01453_),
    .Y(_01674_)
  );
  NAND _09821_ (
    .A(\memory[13][2] ),
    .B(_01520_),
    .Y(_01675_)
  );
  AND _09822_ (
    .A(_01674_),
    .B(_01675_),
    .Y(_01676_)
  );
  AND _09823_ (
    .A(_01673_),
    .B(_01676_),
    .Y(_01677_)
  );
  NAND _09824_ (
    .A(\memory[8][2] ),
    .B(_01527_),
    .Y(_01678_)
  );
  NAND _09825_ (
    .A(\memory[14][2] ),
    .B(_01543_),
    .Y(_01679_)
  );
  AND _09826_ (
    .A(_01678_),
    .B(_01679_),
    .Y(_01680_)
  );
  NAND _09827_ (
    .A(\memory[30][2] ),
    .B(_01491_),
    .Y(_01681_)
  );
  NAND _09828_ (
    .A(\memory[24][2] ),
    .B(_01550_),
    .Y(_01682_)
  );
  AND _09829_ (
    .A(_01681_),
    .B(_01682_),
    .Y(_01683_)
  );
  AND _09830_ (
    .A(_01680_),
    .B(_01683_),
    .Y(_01684_)
  );
  AND _09831_ (
    .A(_01677_),
    .B(_01684_),
    .Y(_01685_)
  );
  AND _09832_ (
    .A(_01670_),
    .B(_01685_),
    .Y(_01686_)
  );
  NAND _09833_ (
    .A(\memory[12][2] ),
    .B(_01458_),
    .Y(_01687_)
  );
  NAND _09834_ (
    .A(\memory[10][2] ),
    .B(_01578_),
    .Y(_01688_)
  );
  AND _09835_ (
    .A(_01687_),
    .B(_01688_),
    .Y(_01689_)
  );
  NAND _09836_ (
    .A(\memory[31][2] ),
    .B(_01504_),
    .Y(_01690_)
  );
  NAND _09837_ (
    .A(\memory[23][2] ),
    .B(_01546_),
    .Y(_01691_)
  );
  AND _09838_ (
    .A(_01690_),
    .B(_01691_),
    .Y(_01692_)
  );
  AND _09839_ (
    .A(_01689_),
    .B(_01692_),
    .Y(_01693_)
  );
  NAND _09840_ (
    .A(\memory[27][2] ),
    .B(_01563_),
    .Y(_01694_)
  );
  NAND _09841_ (
    .A(\memory[20][2] ),
    .B(_01553_),
    .Y(_01695_)
  );
  AND _09842_ (
    .A(_01694_),
    .B(_01695_),
    .Y(_01696_)
  );
  NAND _09843_ (
    .A(\memory[25][2] ),
    .B(_01559_),
    .Y(_01697_)
  );
  NAND _09844_ (
    .A(\memory[17][2] ),
    .B(_01479_),
    .Y(_01698_)
  );
  AND _09845_ (
    .A(_01697_),
    .B(_01698_),
    .Y(_01699_)
  );
  AND _09846_ (
    .A(_01696_),
    .B(_01699_),
    .Y(_01700_)
  );
  AND _09847_ (
    .A(_01693_),
    .B(_01700_),
    .Y(_01701_)
  );
  NAND _09848_ (
    .A(\memory[5][2] ),
    .B(_01585_),
    .Y(_01702_)
  );
  NAND _09849_ (
    .A(\memory[1][2] ),
    .B(_01570_),
    .Y(_01703_)
  );
  AND _09850_ (
    .A(_01702_),
    .B(_01703_),
    .Y(_01704_)
  );
  NAND _09851_ (
    .A(\memory[6][2] ),
    .B(_01517_),
    .Y(_01705_)
  );
  NAND _09852_ (
    .A(\memory[3][2] ),
    .B(_01513_),
    .Y(_01706_)
  );
  AND _09853_ (
    .A(_01705_),
    .B(_01706_),
    .Y(_01707_)
  );
  AND _09854_ (
    .A(_01704_),
    .B(_01707_),
    .Y(_01708_)
  );
  NAND _09855_ (
    .A(\memory[18][2] ),
    .B(_01582_),
    .Y(_01709_)
  );
  NAND _09856_ (
    .A(\memory[22][2] ),
    .B(_01469_),
    .Y(_01710_)
  );
  AND _09857_ (
    .A(_01709_),
    .B(_01710_),
    .Y(_01711_)
  );
  NAND _09858_ (
    .A(\memory[16][2] ),
    .B(_01567_),
    .Y(_01712_)
  );
  NAND _09859_ (
    .A(\memory[21][2] ),
    .B(_01474_),
    .Y(_01713_)
  );
  AND _09860_ (
    .A(_01712_),
    .B(_01713_),
    .Y(_01714_)
  );
  AND _09861_ (
    .A(_01711_),
    .B(_01714_),
    .Y(_01715_)
  );
  AND _09862_ (
    .A(_01708_),
    .B(_01715_),
    .Y(_01716_)
  );
  AND _09863_ (
    .A(_01701_),
    .B(_01716_),
    .Y(_01717_)
  );
  NAND _09864_ (
    .A(_01686_),
    .B(_01717_),
    .Y(_01718_)
  );
  AND _09865_ (
    .A(MemRead_i),
    .B(_01718_),
    .Y(\data_o[2] )
  );
  NAND _09866_ (
    .A(\memory[28][3] ),
    .B(_01462_),
    .Y(_01719_)
  );
  NAND _09867_ (
    .A(\memory[17][3] ),
    .B(_01479_),
    .Y(_01720_)
  );
  AND _09868_ (
    .A(_01719_),
    .B(_01720_),
    .Y(_01721_)
  );
  NAND _09869_ (
    .A(\memory[13][3] ),
    .B(_01520_),
    .Y(_01722_)
  );
  NAND _09870_ (
    .A(\memory[12][3] ),
    .B(_01458_),
    .Y(_01723_)
  );
  AND _09871_ (
    .A(_01722_),
    .B(_01723_),
    .Y(_01724_)
  );
  AND _09872_ (
    .A(_01721_),
    .B(_01724_),
    .Y(_01725_)
  );
  NAND _09873_ (
    .A(\memory[11][3] ),
    .B(_01575_),
    .Y(_01726_)
  );
  NAND _09874_ (
    .A(\memory[29][3] ),
    .B(_01510_),
    .Y(_01727_)
  );
  AND _09875_ (
    .A(_01726_),
    .B(_01727_),
    .Y(_01728_)
  );
  NAND _09876_ (
    .A(\memory[0][3] ),
    .B(_01449_),
    .Y(_01729_)
  );
  NAND _09877_ (
    .A(\memory[4][3] ),
    .B(_01530_),
    .Y(_01730_)
  );
  AND _09878_ (
    .A(_01729_),
    .B(_01730_),
    .Y(_01731_)
  );
  AND _09879_ (
    .A(_01728_),
    .B(_01731_),
    .Y(_01732_)
  );
  AND _09880_ (
    .A(_01725_),
    .B(_01732_),
    .Y(_01733_)
  );
  NAND _09881_ (
    .A(\memory[9][3] ),
    .B(_01495_),
    .Y(_01734_)
  );
  NAND _09882_ (
    .A(\memory[27][3] ),
    .B(_01563_),
    .Y(_01735_)
  );
  AND _09883_ (
    .A(_01734_),
    .B(_01735_),
    .Y(_01736_)
  );
  NAND _09884_ (
    .A(\memory[25][3] ),
    .B(_01559_),
    .Y(_01737_)
  );
  NAND _09885_ (
    .A(\memory[31][3] ),
    .B(_01504_),
    .Y(_01738_)
  );
  AND _09886_ (
    .A(_01737_),
    .B(_01738_),
    .Y(_01739_)
  );
  AND _09887_ (
    .A(_01736_),
    .B(_01739_),
    .Y(_01740_)
  );
  NAND _09888_ (
    .A(\memory[30][3] ),
    .B(_01491_),
    .Y(_01741_)
  );
  NAND _09889_ (
    .A(\memory[10][3] ),
    .B(_01578_),
    .Y(_01742_)
  );
  AND _09890_ (
    .A(_01741_),
    .B(_01742_),
    .Y(_01743_)
  );
  NAND _09891_ (
    .A(\memory[16][3] ),
    .B(_01567_),
    .Y(_01744_)
  );
  NAND _09892_ (
    .A(\memory[6][3] ),
    .B(_01517_),
    .Y(_01745_)
  );
  AND _09893_ (
    .A(_01744_),
    .B(_01745_),
    .Y(_01746_)
  );
  AND _09894_ (
    .A(_01743_),
    .B(_01746_),
    .Y(_01747_)
  );
  AND _09895_ (
    .A(_01740_),
    .B(_01747_),
    .Y(_01748_)
  );
  AND _09896_ (
    .A(_01733_),
    .B(_01748_),
    .Y(_01749_)
  );
  NAND _09897_ (
    .A(\memory[15][3] ),
    .B(_01501_),
    .Y(_01750_)
  );
  NAND _09898_ (
    .A(\memory[1][3] ),
    .B(_01570_),
    .Y(_01751_)
  );
  AND _09899_ (
    .A(_01750_),
    .B(_01751_),
    .Y(_01752_)
  );
  NAND _09900_ (
    .A(\memory[23][3] ),
    .B(_01546_),
    .Y(_01753_)
  );
  NAND _09901_ (
    .A(\memory[21][3] ),
    .B(_01474_),
    .Y(_01754_)
  );
  AND _09902_ (
    .A(_01753_),
    .B(_01754_),
    .Y(_01755_)
  );
  AND _09903_ (
    .A(_01752_),
    .B(_01755_),
    .Y(_01756_)
  );
  NAND _09904_ (
    .A(\memory[5][3] ),
    .B(_01585_),
    .Y(_01757_)
  );
  NAND _09905_ (
    .A(\memory[8][3] ),
    .B(_01527_),
    .Y(_01758_)
  );
  AND _09906_ (
    .A(_01757_),
    .B(_01758_),
    .Y(_01759_)
  );
  NAND _09907_ (
    .A(\memory[19][3] ),
    .B(_01534_),
    .Y(_01760_)
  );
  NAND _09908_ (
    .A(\memory[2][3] ),
    .B(_01453_),
    .Y(_01761_)
  );
  AND _09909_ (
    .A(_01760_),
    .B(_01761_),
    .Y(_01762_)
  );
  AND _09910_ (
    .A(_01759_),
    .B(_01762_),
    .Y(_01763_)
  );
  AND _09911_ (
    .A(_01756_),
    .B(_01763_),
    .Y(_01764_)
  );
  NAND _09912_ (
    .A(\memory[14][3] ),
    .B(_01543_),
    .Y(_01765_)
  );
  NAND _09913_ (
    .A(\memory[7][3] ),
    .B(_01538_),
    .Y(_01766_)
  );
  AND _09914_ (
    .A(_01765_),
    .B(_01766_),
    .Y(_01767_)
  );
  NAND _09915_ (
    .A(\memory[3][3] ),
    .B(_01513_),
    .Y(_01768_)
  );
  NAND _09916_ (
    .A(\memory[18][3] ),
    .B(_01582_),
    .Y(_01769_)
  );
  AND _09917_ (
    .A(_01768_),
    .B(_01769_),
    .Y(_01770_)
  );
  AND _09918_ (
    .A(_01767_),
    .B(_01770_),
    .Y(_01771_)
  );
  NAND _09919_ (
    .A(\memory[20][3] ),
    .B(_01553_),
    .Y(_01772_)
  );
  NAND _09920_ (
    .A(\memory[26][3] ),
    .B(_01484_),
    .Y(_01773_)
  );
  AND _09921_ (
    .A(_01772_),
    .B(_01773_),
    .Y(_01774_)
  );
  NAND _09922_ (
    .A(\memory[24][3] ),
    .B(_01550_),
    .Y(_01775_)
  );
  NAND _09923_ (
    .A(\memory[22][3] ),
    .B(_01469_),
    .Y(_01776_)
  );
  AND _09924_ (
    .A(_01775_),
    .B(_01776_),
    .Y(_01777_)
  );
  AND _09925_ (
    .A(_01774_),
    .B(_01777_),
    .Y(_01778_)
  );
  AND _09926_ (
    .A(_01771_),
    .B(_01778_),
    .Y(_01779_)
  );
  AND _09927_ (
    .A(_01764_),
    .B(_01779_),
    .Y(_01780_)
  );
  NAND _09928_ (
    .A(_01749_),
    .B(_01780_),
    .Y(_01781_)
  );
  AND _09929_ (
    .A(MemRead_i),
    .B(_01781_),
    .Y(\data_o[3] )
  );
  NAND _09930_ (
    .A(\memory[28][4] ),
    .B(_01462_),
    .Y(_01782_)
  );
  NAND _09931_ (
    .A(\memory[18][4] ),
    .B(_01582_),
    .Y(_01783_)
  );
  AND _09932_ (
    .A(_01782_),
    .B(_01783_),
    .Y(_01784_)
  );
  NAND _09933_ (
    .A(\memory[20][4] ),
    .B(_01553_),
    .Y(_01785_)
  );
  NAND _09934_ (
    .A(\memory[5][4] ),
    .B(_01585_),
    .Y(_01786_)
  );
  AND _09935_ (
    .A(_01785_),
    .B(_01786_),
    .Y(_01787_)
  );
  AND _09936_ (
    .A(_01784_),
    .B(_01787_),
    .Y(_01788_)
  );
  NAND _09937_ (
    .A(\memory[15][4] ),
    .B(_01501_),
    .Y(_01789_)
  );
  NAND _09938_ (
    .A(\memory[29][4] ),
    .B(_01510_),
    .Y(_01790_)
  );
  AND _09939_ (
    .A(_01789_),
    .B(_01790_),
    .Y(_01791_)
  );
  NAND _09940_ (
    .A(\memory[0][4] ),
    .B(_01449_),
    .Y(_01792_)
  );
  NAND _09941_ (
    .A(\memory[6][4] ),
    .B(_01517_),
    .Y(_01793_)
  );
  AND _09942_ (
    .A(_01792_),
    .B(_01793_),
    .Y(_01794_)
  );
  AND _09943_ (
    .A(_01791_),
    .B(_01794_),
    .Y(_01795_)
  );
  AND _09944_ (
    .A(_01788_),
    .B(_01795_),
    .Y(_01796_)
  );
  NAND _09945_ (
    .A(\memory[13][4] ),
    .B(_01520_),
    .Y(_01797_)
  );
  NAND _09946_ (
    .A(\memory[27][4] ),
    .B(_01563_),
    .Y(_01798_)
  );
  AND _09947_ (
    .A(_01797_),
    .B(_01798_),
    .Y(_01799_)
  );
  NAND _09948_ (
    .A(\memory[25][4] ),
    .B(_01559_),
    .Y(_01800_)
  );
  NAND _09949_ (
    .A(\memory[31][4] ),
    .B(_01504_),
    .Y(_01801_)
  );
  AND _09950_ (
    .A(_01800_),
    .B(_01801_),
    .Y(_01802_)
  );
  AND _09951_ (
    .A(_01799_),
    .B(_01802_),
    .Y(_01803_)
  );
  NAND _09952_ (
    .A(\memory[1][4] ),
    .B(_01570_),
    .Y(_01804_)
  );
  NAND _09953_ (
    .A(\memory[30][4] ),
    .B(_01491_),
    .Y(_01805_)
  );
  AND _09954_ (
    .A(_01804_),
    .B(_01805_),
    .Y(_01806_)
  );
  NAND _09955_ (
    .A(\memory[22][4] ),
    .B(_01469_),
    .Y(_01807_)
  );
  NAND _09956_ (
    .A(\memory[14][4] ),
    .B(_01543_),
    .Y(_01808_)
  );
  AND _09957_ (
    .A(_01807_),
    .B(_01808_),
    .Y(_01809_)
  );
  AND _09958_ (
    .A(_01806_),
    .B(_01809_),
    .Y(_01810_)
  );
  AND _09959_ (
    .A(_01803_),
    .B(_01810_),
    .Y(_01811_)
  );
  AND _09960_ (
    .A(_01796_),
    .B(_01811_),
    .Y(_01812_)
  );
  NAND _09961_ (
    .A(\memory[7][4] ),
    .B(_01538_),
    .Y(_01813_)
  );
  NAND _09962_ (
    .A(\memory[24][4] ),
    .B(_01550_),
    .Y(_01814_)
  );
  AND _09963_ (
    .A(_01813_),
    .B(_01814_),
    .Y(_01815_)
  );
  NAND _09964_ (
    .A(\memory[16][4] ),
    .B(_01567_),
    .Y(_01816_)
  );
  NAND _09965_ (
    .A(\memory[11][4] ),
    .B(_01575_),
    .Y(_01817_)
  );
  AND _09966_ (
    .A(_01816_),
    .B(_01817_),
    .Y(_01818_)
  );
  AND _09967_ (
    .A(_01815_),
    .B(_01818_),
    .Y(_01819_)
  );
  NAND _09968_ (
    .A(\memory[9][4] ),
    .B(_01495_),
    .Y(_01820_)
  );
  NAND _09969_ (
    .A(\memory[19][4] ),
    .B(_01534_),
    .Y(_01821_)
  );
  AND _09970_ (
    .A(_01820_),
    .B(_01821_),
    .Y(_01822_)
  );
  NAND _09971_ (
    .A(\memory[2][4] ),
    .B(_01453_),
    .Y(_01823_)
  );
  NAND _09972_ (
    .A(\memory[21][4] ),
    .B(_01474_),
    .Y(_01824_)
  );
  AND _09973_ (
    .A(_01823_),
    .B(_01824_),
    .Y(_01825_)
  );
  AND _09974_ (
    .A(_01822_),
    .B(_01825_),
    .Y(_01826_)
  );
  AND _09975_ (
    .A(_01819_),
    .B(_01826_),
    .Y(_01827_)
  );
  NAND _09976_ (
    .A(\memory[23][4] ),
    .B(_01546_),
    .Y(_01828_)
  );
  NAND _09977_ (
    .A(\memory[10][4] ),
    .B(_01578_),
    .Y(_01829_)
  );
  AND _09978_ (
    .A(_01828_),
    .B(_01829_),
    .Y(_01830_)
  );
  NAND _09979_ (
    .A(\memory[3][4] ),
    .B(_01513_),
    .Y(_01831_)
  );
  NAND _09980_ (
    .A(\memory[17][4] ),
    .B(_01479_),
    .Y(_01832_)
  );
  AND _09981_ (
    .A(_01831_),
    .B(_01832_),
    .Y(_01833_)
  );
  AND _09982_ (
    .A(_01830_),
    .B(_01833_),
    .Y(_01834_)
  );
  NAND _09983_ (
    .A(\memory[12][4] ),
    .B(_01458_),
    .Y(_01835_)
  );
  NAND _09984_ (
    .A(\memory[4][4] ),
    .B(_01530_),
    .Y(_01836_)
  );
  AND _09985_ (
    .A(_01835_),
    .B(_01836_),
    .Y(_01837_)
  );
  NAND _09986_ (
    .A(\memory[8][4] ),
    .B(_01527_),
    .Y(_01838_)
  );
  NAND _09987_ (
    .A(\memory[26][4] ),
    .B(_01484_),
    .Y(_01839_)
  );
  AND _09988_ (
    .A(_01838_),
    .B(_01839_),
    .Y(_01840_)
  );
  AND _09989_ (
    .A(_01837_),
    .B(_01840_),
    .Y(_01841_)
  );
  AND _09990_ (
    .A(_01834_),
    .B(_01841_),
    .Y(_01842_)
  );
  AND _09991_ (
    .A(_01827_),
    .B(_01842_),
    .Y(_01843_)
  );
  NAND _09992_ (
    .A(_01812_),
    .B(_01843_),
    .Y(_01844_)
  );
  AND _09993_ (
    .A(MemRead_i),
    .B(_01844_),
    .Y(\data_o[4] )
  );
  NAND _09994_ (
    .A(\memory[29][5] ),
    .B(_01510_),
    .Y(_01845_)
  );
  NAND _09995_ (
    .A(\memory[3][5] ),
    .B(_01513_),
    .Y(_01846_)
  );
  AND _09996_ (
    .A(_01845_),
    .B(_01846_),
    .Y(_01847_)
  );
  NAND _09997_ (
    .A(\memory[10][5] ),
    .B(_01578_),
    .Y(_01848_)
  );
  NAND _09998_ (
    .A(\memory[9][5] ),
    .B(_01495_),
    .Y(_01849_)
  );
  AND _09999_ (
    .A(_01848_),
    .B(_01849_),
    .Y(_01850_)
  );
  AND _10000_ (
    .A(_01847_),
    .B(_01850_),
    .Y(_01851_)
  );
  NAND _10001_ (
    .A(\memory[2][5] ),
    .B(_01453_),
    .Y(_01852_)
  );
  NAND _10002_ (
    .A(\memory[6][5] ),
    .B(_01517_),
    .Y(_01853_)
  );
  AND _10003_ (
    .A(_01852_),
    .B(_01853_),
    .Y(_01854_)
  );
  NAND _10004_ (
    .A(\memory[28][5] ),
    .B(_01462_),
    .Y(_01855_)
  );
  NAND _10005_ (
    .A(\memory[0][5] ),
    .B(_01449_),
    .Y(_01856_)
  );
  AND _10006_ (
    .A(_01855_),
    .B(_01856_),
    .Y(_01857_)
  );
  AND _10007_ (
    .A(_01854_),
    .B(_01857_),
    .Y(_01858_)
  );
  AND _10008_ (
    .A(_01851_),
    .B(_01858_),
    .Y(_01859_)
  );
  NAND _10009_ (
    .A(\memory[15][5] ),
    .B(_01501_),
    .Y(_01860_)
  );
  NAND _10010_ (
    .A(\memory[26][5] ),
    .B(_01484_),
    .Y(_01861_)
  );
  AND _10011_ (
    .A(_01860_),
    .B(_01861_),
    .Y(_01862_)
  );
  NAND _10012_ (
    .A(\memory[4][5] ),
    .B(_01530_),
    .Y(_01863_)
  );
  NAND _10013_ (
    .A(\memory[13][5] ),
    .B(_01520_),
    .Y(_01864_)
  );
  AND _10014_ (
    .A(_01863_),
    .B(_01864_),
    .Y(_01865_)
  );
  AND _10015_ (
    .A(_01862_),
    .B(_01865_),
    .Y(_01866_)
  );
  NAND _10016_ (
    .A(\memory[7][5] ),
    .B(_01538_),
    .Y(_01867_)
  );
  NAND _10017_ (
    .A(\memory[14][5] ),
    .B(_01543_),
    .Y(_01868_)
  );
  AND _10018_ (
    .A(_01867_),
    .B(_01868_),
    .Y(_01869_)
  );
  NAND _10019_ (
    .A(\memory[30][5] ),
    .B(_01491_),
    .Y(_01870_)
  );
  NAND _10020_ (
    .A(\memory[24][5] ),
    .B(_01550_),
    .Y(_01871_)
  );
  AND _10021_ (
    .A(_01870_),
    .B(_01871_),
    .Y(_01872_)
  );
  AND _10022_ (
    .A(_01869_),
    .B(_01872_),
    .Y(_01873_)
  );
  AND _10023_ (
    .A(_01866_),
    .B(_01873_),
    .Y(_01874_)
  );
  AND _10024_ (
    .A(_01859_),
    .B(_01874_),
    .Y(_01875_)
  );
  NAND _10025_ (
    .A(\memory[12][5] ),
    .B(_01458_),
    .Y(_01876_)
  );
  NAND _10026_ (
    .A(\memory[16][5] ),
    .B(_01567_),
    .Y(_01877_)
  );
  AND _10027_ (
    .A(_01876_),
    .B(_01877_),
    .Y(_01878_)
  );
  NAND _10028_ (
    .A(\memory[31][5] ),
    .B(_01504_),
    .Y(_01879_)
  );
  NAND _10029_ (
    .A(\memory[23][5] ),
    .B(_01546_),
    .Y(_01880_)
  );
  AND _10030_ (
    .A(_01879_),
    .B(_01880_),
    .Y(_01881_)
  );
  AND _10031_ (
    .A(_01878_),
    .B(_01881_),
    .Y(_01882_)
  );
  NAND _10032_ (
    .A(\memory[27][5] ),
    .B(_01563_),
    .Y(_01883_)
  );
  NAND _10033_ (
    .A(\memory[19][5] ),
    .B(_01534_),
    .Y(_01884_)
  );
  AND _10034_ (
    .A(_01883_),
    .B(_01884_),
    .Y(_01885_)
  );
  NAND _10035_ (
    .A(\memory[25][5] ),
    .B(_01559_),
    .Y(_01886_)
  );
  NAND _10036_ (
    .A(\memory[17][5] ),
    .B(_01479_),
    .Y(_01887_)
  );
  AND _10037_ (
    .A(_01886_),
    .B(_01887_),
    .Y(_01888_)
  );
  AND _10038_ (
    .A(_01885_),
    .B(_01888_),
    .Y(_01889_)
  );
  AND _10039_ (
    .A(_01882_),
    .B(_01889_),
    .Y(_01890_)
  );
  NAND _10040_ (
    .A(\memory[5][5] ),
    .B(_01585_),
    .Y(_01891_)
  );
  NAND _10041_ (
    .A(\memory[8][5] ),
    .B(_01527_),
    .Y(_01892_)
  );
  AND _10042_ (
    .A(_01891_),
    .B(_01892_),
    .Y(_01893_)
  );
  NAND _10043_ (
    .A(\memory[20][5] ),
    .B(_01553_),
    .Y(_01894_)
  );
  NAND _10044_ (
    .A(\memory[1][5] ),
    .B(_01570_),
    .Y(_01895_)
  );
  AND _10045_ (
    .A(_01894_),
    .B(_01895_),
    .Y(_01896_)
  );
  AND _10046_ (
    .A(_01893_),
    .B(_01896_),
    .Y(_01897_)
  );
  NAND _10047_ (
    .A(\memory[18][5] ),
    .B(_01582_),
    .Y(_01898_)
  );
  NAND _10048_ (
    .A(\memory[22][5] ),
    .B(_01469_),
    .Y(_01899_)
  );
  AND _10049_ (
    .A(_01898_),
    .B(_01899_),
    .Y(_01900_)
  );
  NAND _10050_ (
    .A(\memory[11][5] ),
    .B(_01575_),
    .Y(_01901_)
  );
  NAND _10051_ (
    .A(\memory[21][5] ),
    .B(_01474_),
    .Y(_01902_)
  );
  AND _10052_ (
    .A(_01901_),
    .B(_01902_),
    .Y(_01903_)
  );
  AND _10053_ (
    .A(_01900_),
    .B(_01903_),
    .Y(_01904_)
  );
  AND _10054_ (
    .A(_01897_),
    .B(_01904_),
    .Y(_01905_)
  );
  AND _10055_ (
    .A(_01890_),
    .B(_01905_),
    .Y(_01906_)
  );
  NAND _10056_ (
    .A(_01875_),
    .B(_01906_),
    .Y(_01907_)
  );
  AND _10057_ (
    .A(MemRead_i),
    .B(_01907_),
    .Y(\data_o[5] )
  );
  NAND _10058_ (
    .A(\memory[0][6] ),
    .B(_01449_),
    .Y(_01908_)
  );
  NAND _10059_ (
    .A(\memory[29][6] ),
    .B(_01510_),
    .Y(_01909_)
  );
  AND _10060_ (
    .A(_01908_),
    .B(_01909_),
    .Y(_01910_)
  );
  NAND _10061_ (
    .A(\memory[31][6] ),
    .B(_01504_),
    .Y(_01911_)
  );
  NAND _10062_ (
    .A(\memory[6][6] ),
    .B(_01517_),
    .Y(_01912_)
  );
  AND _10063_ (
    .A(_01911_),
    .B(_01912_),
    .Y(_01913_)
  );
  AND _10064_ (
    .A(_01910_),
    .B(_01913_),
    .Y(_01914_)
  );
  NAND _10065_ (
    .A(\memory[27][6] ),
    .B(_01563_),
    .Y(_01915_)
  );
  NAND _10066_ (
    .A(\memory[21][6] ),
    .B(_01474_),
    .Y(_01916_)
  );
  AND _10067_ (
    .A(_01915_),
    .B(_01916_),
    .Y(_01917_)
  );
  NAND _10068_ (
    .A(\memory[25][6] ),
    .B(_01559_),
    .Y(_01918_)
  );
  NAND _10069_ (
    .A(\memory[14][6] ),
    .B(_01543_),
    .Y(_01919_)
  );
  AND _10070_ (
    .A(_01918_),
    .B(_01919_),
    .Y(_01920_)
  );
  AND _10071_ (
    .A(_01917_),
    .B(_01920_),
    .Y(_01921_)
  );
  AND _10072_ (
    .A(_01914_),
    .B(_01921_),
    .Y(_01922_)
  );
  NAND _10073_ (
    .A(\memory[8][6] ),
    .B(_01527_),
    .Y(_01923_)
  );
  NAND _10074_ (
    .A(\memory[20][6] ),
    .B(_01553_),
    .Y(_01924_)
  );
  AND _10075_ (
    .A(_01923_),
    .B(_01924_),
    .Y(_01925_)
  );
  NAND _10076_ (
    .A(\memory[19][6] ),
    .B(_01534_),
    .Y(_01926_)
  );
  NAND _10077_ (
    .A(\memory[17][6] ),
    .B(_01479_),
    .Y(_01927_)
  );
  AND _10078_ (
    .A(_01926_),
    .B(_01927_),
    .Y(_01928_)
  );
  AND _10079_ (
    .A(_01925_),
    .B(_01928_),
    .Y(_01929_)
  );
  NAND _10080_ (
    .A(\memory[3][6] ),
    .B(_01513_),
    .Y(_01930_)
  );
  NAND _10081_ (
    .A(\memory[18][6] ),
    .B(_01582_),
    .Y(_01931_)
  );
  AND _10082_ (
    .A(_01930_),
    .B(_01931_),
    .Y(_01932_)
  );
  NAND _10083_ (
    .A(\memory[7][6] ),
    .B(_01538_),
    .Y(_01933_)
  );
  NAND _10084_ (
    .A(\memory[28][6] ),
    .B(_01462_),
    .Y(_01934_)
  );
  AND _10085_ (
    .A(_01933_),
    .B(_01934_),
    .Y(_01935_)
  );
  AND _10086_ (
    .A(_01932_),
    .B(_01935_),
    .Y(_01936_)
  );
  AND _10087_ (
    .A(_01929_),
    .B(_01936_),
    .Y(_01937_)
  );
  AND _10088_ (
    .A(_01922_),
    .B(_01937_),
    .Y(_01938_)
  );
  NAND _10089_ (
    .A(\memory[24][6] ),
    .B(_01550_),
    .Y(_01939_)
  );
  NAND _10090_ (
    .A(\memory[22][6] ),
    .B(_01469_),
    .Y(_01940_)
  );
  AND _10091_ (
    .A(_01939_),
    .B(_01940_),
    .Y(_01941_)
  );
  NAND _10092_ (
    .A(\memory[1][6] ),
    .B(_01570_),
    .Y(_01942_)
  );
  NAND _10093_ (
    .A(\memory[16][6] ),
    .B(_01567_),
    .Y(_01943_)
  );
  AND _10094_ (
    .A(_01942_),
    .B(_01943_),
    .Y(_01944_)
  );
  AND _10095_ (
    .A(_01941_),
    .B(_01944_),
    .Y(_01945_)
  );
  NAND _10096_ (
    .A(\memory[10][6] ),
    .B(_01578_),
    .Y(_01946_)
  );
  NAND _10097_ (
    .A(\memory[9][6] ),
    .B(_01495_),
    .Y(_01947_)
  );
  AND _10098_ (
    .A(_01946_),
    .B(_01947_),
    .Y(_01948_)
  );
  NAND _10099_ (
    .A(\memory[2][6] ),
    .B(_01453_),
    .Y(_01949_)
  );
  NAND _10100_ (
    .A(\memory[4][6] ),
    .B(_01530_),
    .Y(_01950_)
  );
  AND _10101_ (
    .A(_01949_),
    .B(_01950_),
    .Y(_01951_)
  );
  AND _10102_ (
    .A(_01948_),
    .B(_01951_),
    .Y(_01952_)
  );
  AND _10103_ (
    .A(_01945_),
    .B(_01952_),
    .Y(_01953_)
  );
  NAND _10104_ (
    .A(\memory[15][6] ),
    .B(_01501_),
    .Y(_01954_)
  );
  NAND _10105_ (
    .A(\memory[5][6] ),
    .B(_01585_),
    .Y(_01955_)
  );
  AND _10106_ (
    .A(_01954_),
    .B(_01955_),
    .Y(_01956_)
  );
  NAND _10107_ (
    .A(\memory[23][6] ),
    .B(_01546_),
    .Y(_01957_)
  );
  NAND _10108_ (
    .A(\memory[13][6] ),
    .B(_01520_),
    .Y(_01958_)
  );
  AND _10109_ (
    .A(_01957_),
    .B(_01958_),
    .Y(_01959_)
  );
  AND _10110_ (
    .A(_01956_),
    .B(_01959_),
    .Y(_01960_)
  );
  NAND _10111_ (
    .A(\memory[26][6] ),
    .B(_01484_),
    .Y(_01961_)
  );
  NAND _10112_ (
    .A(\memory[30][6] ),
    .B(_01491_),
    .Y(_01962_)
  );
  AND _10113_ (
    .A(_01961_),
    .B(_01962_),
    .Y(_01963_)
  );
  NAND _10114_ (
    .A(\memory[12][6] ),
    .B(_01458_),
    .Y(_01964_)
  );
  NAND _10115_ (
    .A(\memory[11][6] ),
    .B(_01575_),
    .Y(_01965_)
  );
  AND _10116_ (
    .A(_01964_),
    .B(_01965_),
    .Y(_01966_)
  );
  AND _10117_ (
    .A(_01963_),
    .B(_01966_),
    .Y(_01967_)
  );
  AND _10118_ (
    .A(_01960_),
    .B(_01967_),
    .Y(_01968_)
  );
  AND _10119_ (
    .A(_01953_),
    .B(_01968_),
    .Y(_01969_)
  );
  NAND _10120_ (
    .A(_01938_),
    .B(_01969_),
    .Y(_01970_)
  );
  AND _10121_ (
    .A(MemRead_i),
    .B(_01970_),
    .Y(\data_o[6] )
  );
  NAND _10122_ (
    .A(\memory[16][7] ),
    .B(_01567_),
    .Y(_01971_)
  );
  NAND _10123_ (
    .A(\memory[15][7] ),
    .B(_01501_),
    .Y(_01972_)
  );
  AND _10124_ (
    .A(_01971_),
    .B(_01972_),
    .Y(_01973_)
  );
  NAND _10125_ (
    .A(\memory[11][7] ),
    .B(_01575_),
    .Y(_01974_)
  );
  NAND _10126_ (
    .A(\memory[17][7] ),
    .B(_01479_),
    .Y(_01975_)
  );
  AND _10127_ (
    .A(_01974_),
    .B(_01975_),
    .Y(_01976_)
  );
  AND _10128_ (
    .A(_01973_),
    .B(_01976_),
    .Y(_01977_)
  );
  NAND _10129_ (
    .A(\memory[6][7] ),
    .B(_01517_),
    .Y(_01978_)
  );
  NAND _10130_ (
    .A(\memory[21][7] ),
    .B(_01474_),
    .Y(_01979_)
  );
  AND _10131_ (
    .A(_01978_),
    .B(_01979_),
    .Y(_01980_)
  );
  NAND _10132_ (
    .A(\memory[0][7] ),
    .B(_01449_),
    .Y(_01981_)
  );
  NAND _10133_ (
    .A(\memory[3][7] ),
    .B(_01513_),
    .Y(_01982_)
  );
  AND _10134_ (
    .A(_01981_),
    .B(_01982_),
    .Y(_01983_)
  );
  AND _10135_ (
    .A(_01980_),
    .B(_01983_),
    .Y(_01984_)
  );
  AND _10136_ (
    .A(_01977_),
    .B(_01984_),
    .Y(_01985_)
  );
  NAND _10137_ (
    .A(\memory[14][7] ),
    .B(_01543_),
    .Y(_01986_)
  );
  NAND _10138_ (
    .A(\memory[5][7] ),
    .B(_01585_),
    .Y(_01987_)
  );
  AND _10139_ (
    .A(_01986_),
    .B(_01987_),
    .Y(_01988_)
  );
  NAND _10140_ (
    .A(\memory[24][7] ),
    .B(_01550_),
    .Y(_01989_)
  );
  NAND _10141_ (
    .A(\memory[13][7] ),
    .B(_01520_),
    .Y(_01990_)
  );
  AND _10142_ (
    .A(_01989_),
    .B(_01990_),
    .Y(_01991_)
  );
  AND _10143_ (
    .A(_01988_),
    .B(_01991_),
    .Y(_01992_)
  );
  NAND _10144_ (
    .A(\memory[9][7] ),
    .B(_01495_),
    .Y(_01993_)
  );
  NAND _10145_ (
    .A(\memory[10][7] ),
    .B(_01578_),
    .Y(_01994_)
  );
  AND _10146_ (
    .A(_01993_),
    .B(_01994_),
    .Y(_01995_)
  );
  NAND _10147_ (
    .A(\memory[22][7] ),
    .B(_01469_),
    .Y(_01996_)
  );
  NAND _10148_ (
    .A(\memory[26][7] ),
    .B(_01484_),
    .Y(_01997_)
  );
  AND _10149_ (
    .A(_01996_),
    .B(_01997_),
    .Y(_01998_)
  );
  AND _10150_ (
    .A(_01995_),
    .B(_01998_),
    .Y(_01999_)
  );
  AND _10151_ (
    .A(_01992_),
    .B(_01999_),
    .Y(_02000_)
  );
  AND _10152_ (
    .A(_01985_),
    .B(_02000_),
    .Y(_02001_)
  );
  NAND _10153_ (
    .A(\memory[19][7] ),
    .B(_01534_),
    .Y(_02002_)
  );
  NAND _10154_ (
    .A(\memory[4][7] ),
    .B(_01530_),
    .Y(_02003_)
  );
  AND _10155_ (
    .A(_02002_),
    .B(_02003_),
    .Y(_02004_)
  );
  NAND _10156_ (
    .A(\memory[2][7] ),
    .B(_01453_),
    .Y(_02005_)
  );
  NAND _10157_ (
    .A(\memory[8][7] ),
    .B(_01527_),
    .Y(_02006_)
  );
  AND _10158_ (
    .A(_02005_),
    .B(_02006_),
    .Y(_02007_)
  );
  AND _10159_ (
    .A(_02004_),
    .B(_02007_),
    .Y(_02008_)
  );
  NAND _10160_ (
    .A(\memory[20][7] ),
    .B(_01553_),
    .Y(_02009_)
  );
  NAND _10161_ (
    .A(\memory[1][7] ),
    .B(_01570_),
    .Y(_02010_)
  );
  AND _10162_ (
    .A(_02009_),
    .B(_02010_),
    .Y(_02011_)
  );
  NAND _10163_ (
    .A(\memory[27][7] ),
    .B(_01563_),
    .Y(_02012_)
  );
  NAND _10164_ (
    .A(\memory[12][7] ),
    .B(_01458_),
    .Y(_02013_)
  );
  AND _10165_ (
    .A(_02012_),
    .B(_02013_),
    .Y(_02014_)
  );
  AND _10166_ (
    .A(_02011_),
    .B(_02014_),
    .Y(_02015_)
  );
  AND _10167_ (
    .A(_02008_),
    .B(_02015_),
    .Y(_02016_)
  );
  NAND _10168_ (
    .A(\memory[28][7] ),
    .B(_01462_),
    .Y(_02017_)
  );
  NAND _10169_ (
    .A(\memory[29][7] ),
    .B(_01510_),
    .Y(_02018_)
  );
  AND _10170_ (
    .A(_02017_),
    .B(_02018_),
    .Y(_02019_)
  );
  NAND _10171_ (
    .A(\memory[18][7] ),
    .B(_01582_),
    .Y(_02020_)
  );
  NAND _10172_ (
    .A(\memory[7][7] ),
    .B(_01538_),
    .Y(_02021_)
  );
  AND _10173_ (
    .A(_02020_),
    .B(_02021_),
    .Y(_02022_)
  );
  AND _10174_ (
    .A(_02019_),
    .B(_02022_),
    .Y(_02023_)
  );
  NAND _10175_ (
    .A(\memory[31][7] ),
    .B(_01504_),
    .Y(_02024_)
  );
  NAND _10176_ (
    .A(\memory[30][7] ),
    .B(_01491_),
    .Y(_02025_)
  );
  AND _10177_ (
    .A(_02024_),
    .B(_02025_),
    .Y(_02026_)
  );
  NAND _10178_ (
    .A(\memory[23][7] ),
    .B(_01546_),
    .Y(_02027_)
  );
  NAND _10179_ (
    .A(\memory[25][7] ),
    .B(_01559_),
    .Y(_02028_)
  );
  AND _10180_ (
    .A(_02027_),
    .B(_02028_),
    .Y(_02029_)
  );
  AND _10181_ (
    .A(_02026_),
    .B(_02029_),
    .Y(_02030_)
  );
  AND _10182_ (
    .A(_02023_),
    .B(_02030_),
    .Y(_02031_)
  );
  AND _10183_ (
    .A(_02016_),
    .B(_02031_),
    .Y(_02032_)
  );
  NAND _10184_ (
    .A(_02001_),
    .B(_02032_),
    .Y(_02033_)
  );
  AND _10185_ (
    .A(MemRead_i),
    .B(_02033_),
    .Y(\data_o[7] )
  );
  NAND _10186_ (
    .A(\memory[23][0] ),
    .B(_01469_),
    .Y(_02034_)
  );
  NAND _10187_ (
    .A(\memory[15][0] ),
    .B(_01543_),
    .Y(_02035_)
  );
  AND _10188_ (
    .A(_02034_),
    .B(_02035_),
    .Y(_02036_)
  );
  NAND _10189_ (
    .A(\memory[16][0] ),
    .B(_01501_),
    .Y(_02037_)
  );
  NAND _10190_ (
    .A(\memory[14][0] ),
    .B(_01520_),
    .Y(_02038_)
  );
  AND _10191_ (
    .A(_02037_),
    .B(_02038_),
    .Y(_02039_)
  );
  AND _10192_ (
    .A(_02036_),
    .B(_02039_),
    .Y(_02040_)
  );
  NAND _10193_ (
    .A(\memory[11][0] ),
    .B(_01578_),
    .Y(_02041_)
  );
  NAND _10194_ (
    .A(\memory[22][0] ),
    .B(_01474_),
    .Y(_02042_)
  );
  AND _10195_ (
    .A(_02041_),
    .B(_02042_),
    .Y(_02043_)
  );
  NAND _10196_ (
    .A(\memory[20][0] ),
    .B(_01534_),
    .Y(_02044_)
  );
  NAND _10197_ (
    .A(\memory[4][0] ),
    .B(_01513_),
    .Y(_02045_)
  );
  AND _10198_ (
    .A(_02044_),
    .B(_02045_),
    .Y(_02046_)
  );
  AND _10199_ (
    .A(_02043_),
    .B(_02046_),
    .Y(_02047_)
  );
  AND _10200_ (
    .A(_02040_),
    .B(_02047_),
    .Y(_02048_)
  );
  NAND _10201_ (
    .A(\memory[28][0] ),
    .B(_01563_),
    .Y(_02049_)
  );
  NAND _10202_ (
    .A(\memory[2][0] ),
    .B(_01570_),
    .Y(_02050_)
  );
  AND _10203_ (
    .A(_02049_),
    .B(_02050_),
    .Y(_02051_)
  );
  NAND _10204_ (
    .A(\memory[7][0] ),
    .B(_01517_),
    .Y(_02052_)
  );
  NAND _10205_ (
    .A(\memory[24][0] ),
    .B(_01546_),
    .Y(_02053_)
  );
  AND _10206_ (
    .A(_02052_),
    .B(_02053_),
    .Y(_02054_)
  );
  AND _10207_ (
    .A(_02051_),
    .B(_02054_),
    .Y(_02055_)
  );
  NAND _10208_ (
    .A(\memory[10][0] ),
    .B(_01495_),
    .Y(_02056_)
  );
  NAND _10209_ (
    .A(\memory[12][0] ),
    .B(_01575_),
    .Y(_02057_)
  );
  AND _10210_ (
    .A(_02056_),
    .B(_02057_),
    .Y(_02058_)
  );
  NAND _10211_ (
    .A(\memory[1][0] ),
    .B(_01449_),
    .Y(_02059_)
  );
  NAND _10212_ (
    .A(\memory[3][0] ),
    .B(_01453_),
    .Y(_02060_)
  );
  AND _10213_ (
    .A(_02059_),
    .B(_02060_),
    .Y(_02061_)
  );
  AND _10214_ (
    .A(_02058_),
    .B(_02061_),
    .Y(_02062_)
  );
  AND _10215_ (
    .A(_02055_),
    .B(_02062_),
    .Y(_02063_)
  );
  AND _10216_ (
    .A(_02048_),
    .B(_02063_),
    .Y(_02064_)
  );
  NAND _10217_ (
    .A(\memory[8][0] ),
    .B(_01538_),
    .Y(_02065_)
  );
  NAND _10218_ (
    .A(\memory[27][0] ),
    .B(_01484_),
    .Y(_02066_)
  );
  AND _10219_ (
    .A(_02065_),
    .B(_02066_),
    .Y(_02067_)
  );
  NAND _10220_ (
    .A(\memory[17][0] ),
    .B(_01567_),
    .Y(_02068_)
  );
  NAND _10221_ (
    .A(\memory[6][0] ),
    .B(_01585_),
    .Y(_02069_)
  );
  AND _10222_ (
    .A(_02068_),
    .B(_02069_),
    .Y(_02070_)
  );
  AND _10223_ (
    .A(_02067_),
    .B(_02070_),
    .Y(_02071_)
  );
  NAND _10224_ (
    .A(\memory[30][0] ),
    .B(_01510_),
    .Y(_02072_)
  );
  NAND _10225_ (
    .A(\memory[0][0] ),
    .B(_01504_),
    .Y(_02073_)
  );
  AND _10226_ (
    .A(_02072_),
    .B(_02073_),
    .Y(_02074_)
  );
  NAND _10227_ (
    .A(\memory[13][0] ),
    .B(_01458_),
    .Y(_02075_)
  );
  NAND _10228_ (
    .A(\memory[26][0] ),
    .B(_01559_),
    .Y(_02076_)
  );
  AND _10229_ (
    .A(_02075_),
    .B(_02076_),
    .Y(_02077_)
  );
  AND _10230_ (
    .A(_02074_),
    .B(_02077_),
    .Y(_02078_)
  );
  AND _10231_ (
    .A(_02071_),
    .B(_02078_),
    .Y(_02079_)
  );
  NAND _10232_ (
    .A(\memory[9][0] ),
    .B(_01527_),
    .Y(_02080_)
  );
  NAND _10233_ (
    .A(\memory[5][0] ),
    .B(_01530_),
    .Y(_02081_)
  );
  AND _10234_ (
    .A(_02080_),
    .B(_02081_),
    .Y(_02082_)
  );
  NAND _10235_ (
    .A(\memory[29][0] ),
    .B(_01462_),
    .Y(_02083_)
  );
  NAND _10236_ (
    .A(\memory[25][0] ),
    .B(_01550_),
    .Y(_02084_)
  );
  AND _10237_ (
    .A(_02083_),
    .B(_02084_),
    .Y(_02085_)
  );
  AND _10238_ (
    .A(_02082_),
    .B(_02085_),
    .Y(_02086_)
  );
  NAND _10239_ (
    .A(\memory[19][0] ),
    .B(_01582_),
    .Y(_02087_)
  );
  NAND _10240_ (
    .A(\memory[31][0] ),
    .B(_01491_),
    .Y(_02088_)
  );
  AND _10241_ (
    .A(_02087_),
    .B(_02088_),
    .Y(_02089_)
  );
  NAND _10242_ (
    .A(\memory[21][0] ),
    .B(_01553_),
    .Y(_02090_)
  );
  NAND _10243_ (
    .A(\memory[18][0] ),
    .B(_01479_),
    .Y(_02091_)
  );
  AND _10244_ (
    .A(_02090_),
    .B(_02091_),
    .Y(_02092_)
  );
  AND _10245_ (
    .A(_02089_),
    .B(_02092_),
    .Y(_02093_)
  );
  AND _10246_ (
    .A(_02086_),
    .B(_02093_),
    .Y(_02094_)
  );
  AND _10247_ (
    .A(_02079_),
    .B(_02094_),
    .Y(_02095_)
  );
  NAND _10248_ (
    .A(_02064_),
    .B(_02095_),
    .Y(_02096_)
  );
  AND _10249_ (
    .A(MemRead_i),
    .B(_02096_),
    .Y(\data_o[8] )
  );
  NAND _10250_ (
    .A(\memory[31][1] ),
    .B(_01491_),
    .Y(_02097_)
  );
  NAND _10251_ (
    .A(\memory[1][1] ),
    .B(_01449_),
    .Y(_02098_)
  );
  AND _10252_ (
    .A(_02097_),
    .B(_02098_),
    .Y(_02099_)
  );
  NAND _10253_ (
    .A(\memory[4][1] ),
    .B(_01513_),
    .Y(_02100_)
  );
  NAND _10254_ (
    .A(\memory[22][1] ),
    .B(_01474_),
    .Y(_02101_)
  );
  AND _10255_ (
    .A(_02100_),
    .B(_02101_),
    .Y(_02102_)
  );
  AND _10256_ (
    .A(_02099_),
    .B(_02102_),
    .Y(_02103_)
  );
  NAND _10257_ (
    .A(\memory[5][1] ),
    .B(_01530_),
    .Y(_02104_)
  );
  NAND _10258_ (
    .A(\memory[12][1] ),
    .B(_01575_),
    .Y(_02105_)
  );
  AND _10259_ (
    .A(_02104_),
    .B(_02105_),
    .Y(_02106_)
  );
  NAND _10260_ (
    .A(\memory[20][1] ),
    .B(_01534_),
    .Y(_02107_)
  );
  NAND _10261_ (
    .A(\memory[6][1] ),
    .B(_01585_),
    .Y(_02108_)
  );
  AND _10262_ (
    .A(_02107_),
    .B(_02108_),
    .Y(_02109_)
  );
  AND _10263_ (
    .A(_02106_),
    .B(_02109_),
    .Y(_02110_)
  );
  AND _10264_ (
    .A(_02103_),
    .B(_02110_),
    .Y(_02111_)
  );
  NAND _10265_ (
    .A(\memory[7][1] ),
    .B(_01517_),
    .Y(_02112_)
  );
  NAND _10266_ (
    .A(\memory[2][1] ),
    .B(_01570_),
    .Y(_02113_)
  );
  AND _10267_ (
    .A(_02112_),
    .B(_02113_),
    .Y(_02114_)
  );
  NAND _10268_ (
    .A(\memory[28][1] ),
    .B(_01563_),
    .Y(_02115_)
  );
  NAND _10269_ (
    .A(\memory[18][1] ),
    .B(_01479_),
    .Y(_02116_)
  );
  AND _10270_ (
    .A(_02115_),
    .B(_02116_),
    .Y(_02117_)
  );
  AND _10271_ (
    .A(_02114_),
    .B(_02117_),
    .Y(_02118_)
  );
  NAND _10272_ (
    .A(\memory[17][1] ),
    .B(_01567_),
    .Y(_02119_)
  );
  NAND _10273_ (
    .A(\memory[19][1] ),
    .B(_01582_),
    .Y(_02120_)
  );
  AND _10274_ (
    .A(_02119_),
    .B(_02120_),
    .Y(_02121_)
  );
  NAND _10275_ (
    .A(\memory[16][1] ),
    .B(_01501_),
    .Y(_02122_)
  );
  NAND _10276_ (
    .A(\memory[24][1] ),
    .B(_01546_),
    .Y(_02123_)
  );
  AND _10277_ (
    .A(_02122_),
    .B(_02123_),
    .Y(_02124_)
  );
  AND _10278_ (
    .A(_02121_),
    .B(_02124_),
    .Y(_02125_)
  );
  AND _10279_ (
    .A(_02118_),
    .B(_02125_),
    .Y(_02126_)
  );
  AND _10280_ (
    .A(_02111_),
    .B(_02126_),
    .Y(_02127_)
  );
  NAND _10281_ (
    .A(\memory[13][1] ),
    .B(_01458_),
    .Y(_02128_)
  );
  NAND _10282_ (
    .A(\memory[29][1] ),
    .B(_01462_),
    .Y(_02129_)
  );
  AND _10283_ (
    .A(_02128_),
    .B(_02129_),
    .Y(_02130_)
  );
  NAND _10284_ (
    .A(\memory[8][1] ),
    .B(_01538_),
    .Y(_02131_)
  );
  NAND _10285_ (
    .A(\memory[14][1] ),
    .B(_01520_),
    .Y(_02132_)
  );
  AND _10286_ (
    .A(_02131_),
    .B(_02132_),
    .Y(_02133_)
  );
  AND _10287_ (
    .A(_02130_),
    .B(_02133_),
    .Y(_02134_)
  );
  NAND _10288_ (
    .A(\memory[3][1] ),
    .B(_01453_),
    .Y(_02135_)
  );
  NAND _10289_ (
    .A(\memory[9][1] ),
    .B(_01527_),
    .Y(_02136_)
  );
  AND _10290_ (
    .A(_02135_),
    .B(_02136_),
    .Y(_02137_)
  );
  NAND _10291_ (
    .A(\memory[25][1] ),
    .B(_01550_),
    .Y(_02138_)
  );
  NAND _10292_ (
    .A(\memory[21][1] ),
    .B(_01553_),
    .Y(_02139_)
  );
  AND _10293_ (
    .A(_02138_),
    .B(_02139_),
    .Y(_02140_)
  );
  AND _10294_ (
    .A(_02137_),
    .B(_02140_),
    .Y(_02141_)
  );
  AND _10295_ (
    .A(_02134_),
    .B(_02141_),
    .Y(_02142_)
  );
  NAND _10296_ (
    .A(\memory[10][1] ),
    .B(_01495_),
    .Y(_02143_)
  );
  NAND _10297_ (
    .A(\memory[11][1] ),
    .B(_01578_),
    .Y(_02144_)
  );
  AND _10298_ (
    .A(_02143_),
    .B(_02144_),
    .Y(_02145_)
  );
  NAND _10299_ (
    .A(\memory[23][1] ),
    .B(_01469_),
    .Y(_02146_)
  );
  NAND _10300_ (
    .A(\memory[30][1] ),
    .B(_01510_),
    .Y(_02147_)
  );
  AND _10301_ (
    .A(_02146_),
    .B(_02147_),
    .Y(_02148_)
  );
  AND _10302_ (
    .A(_02145_),
    .B(_02148_),
    .Y(_02149_)
  );
  NAND _10303_ (
    .A(\memory[26][1] ),
    .B(_01559_),
    .Y(_02150_)
  );
  NAND _10304_ (
    .A(\memory[0][1] ),
    .B(_01504_),
    .Y(_02151_)
  );
  AND _10305_ (
    .A(_02150_),
    .B(_02151_),
    .Y(_02152_)
  );
  NAND _10306_ (
    .A(\memory[27][1] ),
    .B(_01484_),
    .Y(_02153_)
  );
  NAND _10307_ (
    .A(\memory[15][1] ),
    .B(_01543_),
    .Y(_02154_)
  );
  AND _10308_ (
    .A(_02153_),
    .B(_02154_),
    .Y(_02155_)
  );
  AND _10309_ (
    .A(_02152_),
    .B(_02155_),
    .Y(_02156_)
  );
  AND _10310_ (
    .A(_02149_),
    .B(_02156_),
    .Y(_02157_)
  );
  AND _10311_ (
    .A(_02142_),
    .B(_02157_),
    .Y(_02158_)
  );
  NAND _10312_ (
    .A(_02127_),
    .B(_02158_),
    .Y(_02159_)
  );
  AND _10313_ (
    .A(MemRead_i),
    .B(_02159_),
    .Y(\data_o[9] )
  );
  NAND _10314_ (
    .A(\memory[23][2] ),
    .B(_01469_),
    .Y(_02160_)
  );
  NAND _10315_ (
    .A(\memory[24][2] ),
    .B(_01546_),
    .Y(_02161_)
  );
  AND _10316_ (
    .A(_02160_),
    .B(_02161_),
    .Y(_02162_)
  );
  NAND _10317_ (
    .A(\memory[11][2] ),
    .B(_01578_),
    .Y(_02163_)
  );
  NAND _10318_ (
    .A(\memory[21][2] ),
    .B(_01553_),
    .Y(_02164_)
  );
  AND _10319_ (
    .A(_02163_),
    .B(_02164_),
    .Y(_02165_)
  );
  AND _10320_ (
    .A(_02162_),
    .B(_02165_),
    .Y(_02166_)
  );
  NAND _10321_ (
    .A(\memory[8][2] ),
    .B(_01538_),
    .Y(_02167_)
  );
  NAND _10322_ (
    .A(\memory[15][2] ),
    .B(_01543_),
    .Y(_02168_)
  );
  AND _10323_ (
    .A(_02167_),
    .B(_02168_),
    .Y(_02169_)
  );
  NAND _10324_ (
    .A(\memory[30][2] ),
    .B(_01510_),
    .Y(_02170_)
  );
  NAND _10325_ (
    .A(\memory[25][2] ),
    .B(_01550_),
    .Y(_02171_)
  );
  AND _10326_ (
    .A(_02170_),
    .B(_02171_),
    .Y(_02172_)
  );
  AND _10327_ (
    .A(_02169_),
    .B(_02172_),
    .Y(_02173_)
  );
  AND _10328_ (
    .A(_02166_),
    .B(_02173_),
    .Y(_02174_)
  );
  NAND _10329_ (
    .A(\memory[31][2] ),
    .B(_01491_),
    .Y(_02175_)
  );
  NAND _10330_ (
    .A(\memory[2][2] ),
    .B(_01570_),
    .Y(_02176_)
  );
  AND _10331_ (
    .A(_02175_),
    .B(_02176_),
    .Y(_02177_)
  );
  NAND _10332_ (
    .A(\memory[7][2] ),
    .B(_01517_),
    .Y(_02178_)
  );
  NAND _10333_ (
    .A(\memory[14][2] ),
    .B(_01520_),
    .Y(_02179_)
  );
  AND _10334_ (
    .A(_02178_),
    .B(_02179_),
    .Y(_02180_)
  );
  AND _10335_ (
    .A(_02177_),
    .B(_02180_),
    .Y(_02181_)
  );
  NAND _10336_ (
    .A(\memory[12][2] ),
    .B(_01575_),
    .Y(_02182_)
  );
  NAND _10337_ (
    .A(\memory[27][2] ),
    .B(_01484_),
    .Y(_02183_)
  );
  AND _10338_ (
    .A(_02182_),
    .B(_02183_),
    .Y(_02184_)
  );
  NAND _10339_ (
    .A(\memory[28][2] ),
    .B(_01563_),
    .Y(_02185_)
  );
  NAND _10340_ (
    .A(\memory[29][2] ),
    .B(_01462_),
    .Y(_02186_)
  );
  AND _10341_ (
    .A(_02185_),
    .B(_02186_),
    .Y(_02187_)
  );
  AND _10342_ (
    .A(_02184_),
    .B(_02187_),
    .Y(_02188_)
  );
  AND _10343_ (
    .A(_02181_),
    .B(_02188_),
    .Y(_02189_)
  );
  AND _10344_ (
    .A(_02174_),
    .B(_02189_),
    .Y(_02190_)
  );
  NAND _10345_ (
    .A(\memory[5][2] ),
    .B(_01530_),
    .Y(_02191_)
  );
  NAND _10346_ (
    .A(\memory[10][2] ),
    .B(_01495_),
    .Y(_02192_)
  );
  AND _10347_ (
    .A(_02191_),
    .B(_02192_),
    .Y(_02193_)
  );
  NAND _10348_ (
    .A(\memory[19][2] ),
    .B(_01582_),
    .Y(_02194_)
  );
  NAND _10349_ (
    .A(\memory[0][2] ),
    .B(_01504_),
    .Y(_02195_)
  );
  AND _10350_ (
    .A(_02194_),
    .B(_02195_),
    .Y(_02196_)
  );
  AND _10351_ (
    .A(_02193_),
    .B(_02196_),
    .Y(_02197_)
  );
  NAND _10352_ (
    .A(\memory[17][2] ),
    .B(_01567_),
    .Y(_02198_)
  );
  NAND _10353_ (
    .A(\memory[9][2] ),
    .B(_01527_),
    .Y(_02199_)
  );
  AND _10354_ (
    .A(_02198_),
    .B(_02199_),
    .Y(_02200_)
  );
  NAND _10355_ (
    .A(\memory[6][2] ),
    .B(_01585_),
    .Y(_02201_)
  );
  NAND _10356_ (
    .A(\memory[26][2] ),
    .B(_01559_),
    .Y(_02202_)
  );
  AND _10357_ (
    .A(_02201_),
    .B(_02202_),
    .Y(_02203_)
  );
  AND _10358_ (
    .A(_02200_),
    .B(_02203_),
    .Y(_02204_)
  );
  AND _10359_ (
    .A(_02197_),
    .B(_02204_),
    .Y(_02205_)
  );
  NAND _10360_ (
    .A(\memory[13][2] ),
    .B(_01458_),
    .Y(_02206_)
  );
  NAND _10361_ (
    .A(\memory[22][2] ),
    .B(_01474_),
    .Y(_02207_)
  );
  AND _10362_ (
    .A(_02206_),
    .B(_02207_),
    .Y(_02208_)
  );
  NAND _10363_ (
    .A(\memory[3][2] ),
    .B(_01453_),
    .Y(_02209_)
  );
  NAND _10364_ (
    .A(\memory[16][2] ),
    .B(_01501_),
    .Y(_02210_)
  );
  AND _10365_ (
    .A(_02209_),
    .B(_02210_),
    .Y(_02211_)
  );
  AND _10366_ (
    .A(_02208_),
    .B(_02211_),
    .Y(_02212_)
  );
  NAND _10367_ (
    .A(\memory[20][2] ),
    .B(_01534_),
    .Y(_02213_)
  );
  NAND _10368_ (
    .A(\memory[18][2] ),
    .B(_01479_),
    .Y(_02214_)
  );
  AND _10369_ (
    .A(_02213_),
    .B(_02214_),
    .Y(_02215_)
  );
  NAND _10370_ (
    .A(\memory[1][2] ),
    .B(_01449_),
    .Y(_02216_)
  );
  NAND _10371_ (
    .A(\memory[4][2] ),
    .B(_01513_),
    .Y(_02217_)
  );
  AND _10372_ (
    .A(_02216_),
    .B(_02217_),
    .Y(_02218_)
  );
  AND _10373_ (
    .A(_02215_),
    .B(_02218_),
    .Y(_02219_)
  );
  AND _10374_ (
    .A(_02212_),
    .B(_02219_),
    .Y(_02220_)
  );
  AND _10375_ (
    .A(_02205_),
    .B(_02220_),
    .Y(_02221_)
  );
  NAND _10376_ (
    .A(_02190_),
    .B(_02221_),
    .Y(_02222_)
  );
  AND _10377_ (
    .A(MemRead_i),
    .B(_02222_),
    .Y(\data_o[10] )
  );
  NAND _10378_ (
    .A(\memory[25][3] ),
    .B(_01550_),
    .Y(_02223_)
  );
  NAND _10379_ (
    .A(\memory[24][3] ),
    .B(_01546_),
    .Y(_02224_)
  );
  AND _10380_ (
    .A(_02223_),
    .B(_02224_),
    .Y(_02225_)
  );
  NAND _10381_ (
    .A(\memory[5][3] ),
    .B(_01530_),
    .Y(_02226_)
  );
  NAND _10382_ (
    .A(\memory[27][3] ),
    .B(_01484_),
    .Y(_02227_)
  );
  AND _10383_ (
    .A(_02226_),
    .B(_02227_),
    .Y(_02228_)
  );
  AND _10384_ (
    .A(_02225_),
    .B(_02228_),
    .Y(_02229_)
  );
  NAND _10385_ (
    .A(\memory[26][3] ),
    .B(_01559_),
    .Y(_02230_)
  );
  NAND _10386_ (
    .A(\memory[0][3] ),
    .B(_01504_),
    .Y(_02231_)
  );
  AND _10387_ (
    .A(_02230_),
    .B(_02231_),
    .Y(_02232_)
  );
  NAND _10388_ (
    .A(\memory[30][3] ),
    .B(_01510_),
    .Y(_02233_)
  );
  NAND _10389_ (
    .A(\memory[18][3] ),
    .B(_01479_),
    .Y(_02234_)
  );
  AND _10390_ (
    .A(_02233_),
    .B(_02234_),
    .Y(_02235_)
  );
  AND _10391_ (
    .A(_02232_),
    .B(_02235_),
    .Y(_02236_)
  );
  AND _10392_ (
    .A(_02229_),
    .B(_02236_),
    .Y(_02237_)
  );
  NAND _10393_ (
    .A(\memory[17][3] ),
    .B(_01567_),
    .Y(_02238_)
  );
  NAND _10394_ (
    .A(\memory[16][3] ),
    .B(_01501_),
    .Y(_02239_)
  );
  AND _10395_ (
    .A(_02238_),
    .B(_02239_),
    .Y(_02240_)
  );
  NAND _10396_ (
    .A(\memory[23][3] ),
    .B(_01469_),
    .Y(_02241_)
  );
  NAND _10397_ (
    .A(\memory[15][3] ),
    .B(_01543_),
    .Y(_02242_)
  );
  AND _10398_ (
    .A(_02241_),
    .B(_02242_),
    .Y(_02243_)
  );
  AND _10399_ (
    .A(_02240_),
    .B(_02243_),
    .Y(_02244_)
  );
  NAND _10400_ (
    .A(\memory[20][3] ),
    .B(_01534_),
    .Y(_02245_)
  );
  NAND _10401_ (
    .A(\memory[14][3] ),
    .B(_01520_),
    .Y(_02246_)
  );
  AND _10402_ (
    .A(_02245_),
    .B(_02246_),
    .Y(_02247_)
  );
  NAND _10403_ (
    .A(\memory[11][3] ),
    .B(_01578_),
    .Y(_02248_)
  );
  NAND _10404_ (
    .A(\memory[10][3] ),
    .B(_01495_),
    .Y(_02249_)
  );
  AND _10405_ (
    .A(_02248_),
    .B(_02249_),
    .Y(_02250_)
  );
  AND _10406_ (
    .A(_02247_),
    .B(_02250_),
    .Y(_02251_)
  );
  AND _10407_ (
    .A(_02244_),
    .B(_02251_),
    .Y(_02252_)
  );
  AND _10408_ (
    .A(_02237_),
    .B(_02252_),
    .Y(_02253_)
  );
  NAND _10409_ (
    .A(\memory[2][3] ),
    .B(_01570_),
    .Y(_02254_)
  );
  NAND _10410_ (
    .A(\memory[9][3] ),
    .B(_01527_),
    .Y(_02255_)
  );
  AND _10411_ (
    .A(_02254_),
    .B(_02255_),
    .Y(_02256_)
  );
  NAND _10412_ (
    .A(\memory[22][3] ),
    .B(_01474_),
    .Y(_02257_)
  );
  NAND _10413_ (
    .A(\memory[1][3] ),
    .B(_01449_),
    .Y(_02258_)
  );
  AND _10414_ (
    .A(_02257_),
    .B(_02258_),
    .Y(_02259_)
  );
  AND _10415_ (
    .A(_02256_),
    .B(_02259_),
    .Y(_02260_)
  );
  NAND _10416_ (
    .A(\memory[8][3] ),
    .B(_01538_),
    .Y(_02261_)
  );
  NAND _10417_ (
    .A(\memory[12][3] ),
    .B(_01575_),
    .Y(_02262_)
  );
  AND _10418_ (
    .A(_02261_),
    .B(_02262_),
    .Y(_02263_)
  );
  NAND _10419_ (
    .A(\memory[3][3] ),
    .B(_01453_),
    .Y(_02264_)
  );
  NAND _10420_ (
    .A(\memory[4][3] ),
    .B(_01513_),
    .Y(_02265_)
  );
  AND _10421_ (
    .A(_02264_),
    .B(_02265_),
    .Y(_02266_)
  );
  AND _10422_ (
    .A(_02263_),
    .B(_02266_),
    .Y(_02267_)
  );
  AND _10423_ (
    .A(_02260_),
    .B(_02267_),
    .Y(_02268_)
  );
  NAND _10424_ (
    .A(\memory[21][3] ),
    .B(_01553_),
    .Y(_02269_)
  );
  NAND _10425_ (
    .A(\memory[29][3] ),
    .B(_01462_),
    .Y(_02270_)
  );
  AND _10426_ (
    .A(_02269_),
    .B(_02270_),
    .Y(_02271_)
  );
  NAND _10427_ (
    .A(\memory[13][3] ),
    .B(_01458_),
    .Y(_02272_)
  );
  NAND _10428_ (
    .A(\memory[31][3] ),
    .B(_01491_),
    .Y(_02273_)
  );
  AND _10429_ (
    .A(_02272_),
    .B(_02273_),
    .Y(_02274_)
  );
  AND _10430_ (
    .A(_02271_),
    .B(_02274_),
    .Y(_02275_)
  );
  NAND _10431_ (
    .A(\memory[19][3] ),
    .B(_01582_),
    .Y(_02276_)
  );
  NAND _10432_ (
    .A(\memory[28][3] ),
    .B(_01563_),
    .Y(_02277_)
  );
  AND _10433_ (
    .A(_02276_),
    .B(_02277_),
    .Y(_02278_)
  );
  NAND _10434_ (
    .A(\memory[6][3] ),
    .B(_01585_),
    .Y(_02279_)
  );
  NAND _10435_ (
    .A(\memory[7][3] ),
    .B(_01517_),
    .Y(_02280_)
  );
  AND _10436_ (
    .A(_02279_),
    .B(_02280_),
    .Y(_02281_)
  );
  AND _10437_ (
    .A(_02278_),
    .B(_02281_),
    .Y(_02282_)
  );
  AND _10438_ (
    .A(_02275_),
    .B(_02282_),
    .Y(_02283_)
  );
  AND _10439_ (
    .A(_02268_),
    .B(_02283_),
    .Y(_02284_)
  );
  NAND _10440_ (
    .A(_02253_),
    .B(_02284_),
    .Y(_02285_)
  );
  AND _10441_ (
    .A(MemRead_i),
    .B(_02285_),
    .Y(\data_o[11] )
  );
  NAND _10442_ (
    .A(\memory[26][4] ),
    .B(_01559_),
    .Y(_02286_)
  );
  NAND _10443_ (
    .A(\memory[8][4] ),
    .B(_01538_),
    .Y(_02287_)
  );
  AND _10444_ (
    .A(_02286_),
    .B(_02287_),
    .Y(_02288_)
  );
  NAND _10445_ (
    .A(\memory[25][4] ),
    .B(_01550_),
    .Y(_02289_)
  );
  NAND _10446_ (
    .A(\memory[24][4] ),
    .B(_01546_),
    .Y(_02290_)
  );
  AND _10447_ (
    .A(_02289_),
    .B(_02290_),
    .Y(_02291_)
  );
  AND _10448_ (
    .A(_02288_),
    .B(_02291_),
    .Y(_02292_)
  );
  NAND _10449_ (
    .A(\memory[22][4] ),
    .B(_01474_),
    .Y(_02293_)
  );
  NAND _10450_ (
    .A(\memory[4][4] ),
    .B(_01513_),
    .Y(_02294_)
  );
  AND _10451_ (
    .A(_02293_),
    .B(_02294_),
    .Y(_02295_)
  );
  NAND _10452_ (
    .A(\memory[2][4] ),
    .B(_01570_),
    .Y(_02296_)
  );
  NAND _10453_ (
    .A(\memory[20][4] ),
    .B(_01534_),
    .Y(_02297_)
  );
  AND _10454_ (
    .A(_02296_),
    .B(_02297_),
    .Y(_02298_)
  );
  AND _10455_ (
    .A(_02295_),
    .B(_02298_),
    .Y(_02299_)
  );
  AND _10456_ (
    .A(_02292_),
    .B(_02299_),
    .Y(_02300_)
  );
  NAND _10457_ (
    .A(\memory[14][4] ),
    .B(_01520_),
    .Y(_02301_)
  );
  NAND _10458_ (
    .A(\memory[17][4] ),
    .B(_01567_),
    .Y(_02302_)
  );
  AND _10459_ (
    .A(_02301_),
    .B(_02302_),
    .Y(_02303_)
  );
  NAND _10460_ (
    .A(\memory[0][4] ),
    .B(_01504_),
    .Y(_02304_)
  );
  NAND _10461_ (
    .A(\memory[28][4] ),
    .B(_01563_),
    .Y(_02305_)
  );
  AND _10462_ (
    .A(_02304_),
    .B(_02305_),
    .Y(_02306_)
  );
  AND _10463_ (
    .A(_02303_),
    .B(_02306_),
    .Y(_02307_)
  );
  NAND _10464_ (
    .A(\memory[23][4] ),
    .B(_01469_),
    .Y(_02308_)
  );
  NAND _10465_ (
    .A(\memory[27][4] ),
    .B(_01484_),
    .Y(_02309_)
  );
  AND _10466_ (
    .A(_02308_),
    .B(_02309_),
    .Y(_02310_)
  );
  NAND _10467_ (
    .A(\memory[5][4] ),
    .B(_01530_),
    .Y(_02311_)
  );
  NAND _10468_ (
    .A(\memory[30][4] ),
    .B(_01510_),
    .Y(_02312_)
  );
  AND _10469_ (
    .A(_02311_),
    .B(_02312_),
    .Y(_02313_)
  );
  AND _10470_ (
    .A(_02310_),
    .B(_02313_),
    .Y(_02314_)
  );
  AND _10471_ (
    .A(_02307_),
    .B(_02314_),
    .Y(_02315_)
  );
  AND _10472_ (
    .A(_02300_),
    .B(_02315_),
    .Y(_02316_)
  );
  NAND _10473_ (
    .A(\memory[7][4] ),
    .B(_01517_),
    .Y(_02317_)
  );
  NAND _10474_ (
    .A(\memory[16][4] ),
    .B(_01501_),
    .Y(_02318_)
  );
  AND _10475_ (
    .A(_02317_),
    .B(_02318_),
    .Y(_02319_)
  );
  NAND _10476_ (
    .A(\memory[13][4] ),
    .B(_01458_),
    .Y(_02320_)
  );
  NAND _10477_ (
    .A(\memory[18][4] ),
    .B(_01479_),
    .Y(_02321_)
  );
  AND _10478_ (
    .A(_02320_),
    .B(_02321_),
    .Y(_02322_)
  );
  AND _10479_ (
    .A(_02319_),
    .B(_02322_),
    .Y(_02323_)
  );
  NAND _10480_ (
    .A(\memory[11][4] ),
    .B(_01578_),
    .Y(_02324_)
  );
  NAND _10481_ (
    .A(\memory[12][4] ),
    .B(_01575_),
    .Y(_02325_)
  );
  AND _10482_ (
    .A(_02324_),
    .B(_02325_),
    .Y(_02326_)
  );
  NAND _10483_ (
    .A(\memory[1][4] ),
    .B(_01449_),
    .Y(_02327_)
  );
  NAND _10484_ (
    .A(\memory[29][4] ),
    .B(_01462_),
    .Y(_02328_)
  );
  AND _10485_ (
    .A(_02327_),
    .B(_02328_),
    .Y(_02329_)
  );
  AND _10486_ (
    .A(_02326_),
    .B(_02329_),
    .Y(_02330_)
  );
  AND _10487_ (
    .A(_02323_),
    .B(_02330_),
    .Y(_02331_)
  );
  NAND _10488_ (
    .A(\memory[6][4] ),
    .B(_01585_),
    .Y(_02332_)
  );
  NAND _10489_ (
    .A(\memory[9][4] ),
    .B(_01527_),
    .Y(_02333_)
  );
  AND _10490_ (
    .A(_02332_),
    .B(_02333_),
    .Y(_02334_)
  );
  NAND _10491_ (
    .A(\memory[3][4] ),
    .B(_01453_),
    .Y(_02335_)
  );
  NAND _10492_ (
    .A(\memory[19][4] ),
    .B(_01582_),
    .Y(_02336_)
  );
  AND _10493_ (
    .A(_02335_),
    .B(_02336_),
    .Y(_02337_)
  );
  AND _10494_ (
    .A(_02334_),
    .B(_02337_),
    .Y(_02338_)
  );
  NAND _10495_ (
    .A(\memory[31][4] ),
    .B(_01491_),
    .Y(_02339_)
  );
  NAND _10496_ (
    .A(\memory[10][4] ),
    .B(_01495_),
    .Y(_02340_)
  );
  AND _10497_ (
    .A(_02339_),
    .B(_02340_),
    .Y(_02341_)
  );
  NAND _10498_ (
    .A(\memory[21][4] ),
    .B(_01553_),
    .Y(_02342_)
  );
  NAND _10499_ (
    .A(\memory[15][4] ),
    .B(_01543_),
    .Y(_02343_)
  );
  AND _10500_ (
    .A(_02342_),
    .B(_02343_),
    .Y(_02344_)
  );
  AND _10501_ (
    .A(_02341_),
    .B(_02344_),
    .Y(_02345_)
  );
  AND _10502_ (
    .A(_02338_),
    .B(_02345_),
    .Y(_02346_)
  );
  AND _10503_ (
    .A(_02331_),
    .B(_02346_),
    .Y(_02347_)
  );
  NAND _10504_ (
    .A(_02316_),
    .B(_02347_),
    .Y(_02348_)
  );
  AND _10505_ (
    .A(MemRead_i),
    .B(_02348_),
    .Y(\data_o[12] )
  );
  NAND _10506_ (
    .A(\memory[7][5] ),
    .B(_01517_),
    .Y(_02349_)
  );
  NAND _10507_ (
    .A(\memory[20][5] ),
    .B(_01534_),
    .Y(_02350_)
  );
  AND _10508_ (
    .A(_02349_),
    .B(_02350_),
    .Y(_02351_)
  );
  NAND _10509_ (
    .A(\memory[21][5] ),
    .B(_01553_),
    .Y(_02352_)
  );
  NAND _10510_ (
    .A(\memory[6][5] ),
    .B(_01585_),
    .Y(_02353_)
  );
  AND _10511_ (
    .A(_02352_),
    .B(_02353_),
    .Y(_02354_)
  );
  AND _10512_ (
    .A(_02351_),
    .B(_02354_),
    .Y(_02355_)
  );
  NAND _10513_ (
    .A(\memory[22][5] ),
    .B(_01474_),
    .Y(_02356_)
  );
  NAND _10514_ (
    .A(\memory[26][5] ),
    .B(_01559_),
    .Y(_02357_)
  );
  AND _10515_ (
    .A(_02356_),
    .B(_02357_),
    .Y(_02358_)
  );
  NAND _10516_ (
    .A(\memory[19][5] ),
    .B(_01582_),
    .Y(_02359_)
  );
  NAND _10517_ (
    .A(\memory[24][5] ),
    .B(_01546_),
    .Y(_02360_)
  );
  AND _10518_ (
    .A(_02359_),
    .B(_02360_),
    .Y(_02361_)
  );
  AND _10519_ (
    .A(_02358_),
    .B(_02361_),
    .Y(_02362_)
  );
  AND _10520_ (
    .A(_02355_),
    .B(_02362_),
    .Y(_02363_)
  );
  NAND _10521_ (
    .A(\memory[2][5] ),
    .B(_01570_),
    .Y(_02364_)
  );
  NAND _10522_ (
    .A(\memory[8][5] ),
    .B(_01538_),
    .Y(_02365_)
  );
  AND _10523_ (
    .A(_02364_),
    .B(_02365_),
    .Y(_02366_)
  );
  NAND _10524_ (
    .A(\memory[1][5] ),
    .B(_01449_),
    .Y(_02367_)
  );
  NAND _10525_ (
    .A(\memory[14][5] ),
    .B(_01520_),
    .Y(_02368_)
  );
  AND _10526_ (
    .A(_02367_),
    .B(_02368_),
    .Y(_02369_)
  );
  AND _10527_ (
    .A(_02366_),
    .B(_02369_),
    .Y(_02370_)
  );
  NAND _10528_ (
    .A(\memory[3][5] ),
    .B(_01453_),
    .Y(_02371_)
  );
  NAND _10529_ (
    .A(\memory[4][5] ),
    .B(_01513_),
    .Y(_02372_)
  );
  AND _10530_ (
    .A(_02371_),
    .B(_02372_),
    .Y(_02373_)
  );
  NAND _10531_ (
    .A(\memory[27][5] ),
    .B(_01484_),
    .Y(_02374_)
  );
  NAND _10532_ (
    .A(\memory[30][5] ),
    .B(_01510_),
    .Y(_02375_)
  );
  AND _10533_ (
    .A(_02374_),
    .B(_02375_),
    .Y(_02376_)
  );
  AND _10534_ (
    .A(_02373_),
    .B(_02376_),
    .Y(_02377_)
  );
  AND _10535_ (
    .A(_02370_),
    .B(_02377_),
    .Y(_02378_)
  );
  AND _10536_ (
    .A(_02363_),
    .B(_02378_),
    .Y(_02379_)
  );
  NAND _10537_ (
    .A(\memory[25][5] ),
    .B(_01550_),
    .Y(_02380_)
  );
  NAND _10538_ (
    .A(\memory[5][5] ),
    .B(_01530_),
    .Y(_02381_)
  );
  AND _10539_ (
    .A(_02380_),
    .B(_02381_),
    .Y(_02382_)
  );
  NAND _10540_ (
    .A(\memory[16][5] ),
    .B(_01501_),
    .Y(_02383_)
  );
  NAND _10541_ (
    .A(\memory[18][5] ),
    .B(_01479_),
    .Y(_02384_)
  );
  AND _10542_ (
    .A(_02383_),
    .B(_02384_),
    .Y(_02385_)
  );
  AND _10543_ (
    .A(_02382_),
    .B(_02385_),
    .Y(_02386_)
  );
  NAND _10544_ (
    .A(\memory[17][5] ),
    .B(_01567_),
    .Y(_02387_)
  );
  NAND _10545_ (
    .A(\memory[28][5] ),
    .B(_01563_),
    .Y(_02388_)
  );
  AND _10546_ (
    .A(_02387_),
    .B(_02388_),
    .Y(_02389_)
  );
  NAND _10547_ (
    .A(\memory[9][5] ),
    .B(_01527_),
    .Y(_02390_)
  );
  NAND _10548_ (
    .A(\memory[31][5] ),
    .B(_01491_),
    .Y(_02391_)
  );
  AND _10549_ (
    .A(_02390_),
    .B(_02391_),
    .Y(_02392_)
  );
  AND _10550_ (
    .A(_02389_),
    .B(_02392_),
    .Y(_02393_)
  );
  AND _10551_ (
    .A(_02386_),
    .B(_02393_),
    .Y(_02394_)
  );
  NAND _10552_ (
    .A(\memory[12][5] ),
    .B(_01575_),
    .Y(_02395_)
  );
  NAND _10553_ (
    .A(\memory[10][5] ),
    .B(_01495_),
    .Y(_02396_)
  );
  AND _10554_ (
    .A(_02395_),
    .B(_02396_),
    .Y(_02397_)
  );
  NAND _10555_ (
    .A(\memory[23][5] ),
    .B(_01469_),
    .Y(_02398_)
  );
  NAND _10556_ (
    .A(\memory[0][5] ),
    .B(_01504_),
    .Y(_02399_)
  );
  AND _10557_ (
    .A(_02398_),
    .B(_02399_),
    .Y(_02400_)
  );
  AND _10558_ (
    .A(_02397_),
    .B(_02400_),
    .Y(_02401_)
  );
  NAND _10559_ (
    .A(\memory[13][5] ),
    .B(_01458_),
    .Y(_02402_)
  );
  NAND _10560_ (
    .A(\memory[15][5] ),
    .B(_01543_),
    .Y(_02403_)
  );
  AND _10561_ (
    .A(_02402_),
    .B(_02403_),
    .Y(_02404_)
  );
  NAND _10562_ (
    .A(\memory[29][5] ),
    .B(_01462_),
    .Y(_02405_)
  );
  NAND _10563_ (
    .A(\memory[11][5] ),
    .B(_01578_),
    .Y(_02406_)
  );
  AND _10564_ (
    .A(_02405_),
    .B(_02406_),
    .Y(_02407_)
  );
  AND _10565_ (
    .A(_02404_),
    .B(_02407_),
    .Y(_02408_)
  );
  AND _10566_ (
    .A(_02401_),
    .B(_02408_),
    .Y(_02409_)
  );
  AND _10567_ (
    .A(_02394_),
    .B(_02409_),
    .Y(_02410_)
  );
  NAND _10568_ (
    .A(_02379_),
    .B(_02410_),
    .Y(_02411_)
  );
  AND _10569_ (
    .A(MemRead_i),
    .B(_02411_),
    .Y(\data_o[13] )
  );
  NAND _10570_ (
    .A(\memory[5][6] ),
    .B(_01530_),
    .Y(_02412_)
  );
  NAND _10571_ (
    .A(\memory[1][6] ),
    .B(_01449_),
    .Y(_02413_)
  );
  AND _10572_ (
    .A(_02412_),
    .B(_02413_),
    .Y(_02414_)
  );
  NAND _10573_ (
    .A(\memory[15][6] ),
    .B(_01543_),
    .Y(_02415_)
  );
  NAND _10574_ (
    .A(\memory[6][6] ),
    .B(_01585_),
    .Y(_02416_)
  );
  AND _10575_ (
    .A(_02415_),
    .B(_02416_),
    .Y(_02417_)
  );
  AND _10576_ (
    .A(_02414_),
    .B(_02417_),
    .Y(_02418_)
  );
  NAND _10577_ (
    .A(\memory[21][6] ),
    .B(_01553_),
    .Y(_02419_)
  );
  NAND _10578_ (
    .A(\memory[0][6] ),
    .B(_01504_),
    .Y(_02420_)
  );
  AND _10579_ (
    .A(_02419_),
    .B(_02420_),
    .Y(_02421_)
  );
  NAND _10580_ (
    .A(\memory[29][6] ),
    .B(_01462_),
    .Y(_02422_)
  );
  NAND _10581_ (
    .A(\memory[30][6] ),
    .B(_01510_),
    .Y(_02423_)
  );
  AND _10582_ (
    .A(_02422_),
    .B(_02423_),
    .Y(_02424_)
  );
  AND _10583_ (
    .A(_02421_),
    .B(_02424_),
    .Y(_02425_)
  );
  AND _10584_ (
    .A(_02418_),
    .B(_02425_),
    .Y(_02426_)
  );
  NAND _10585_ (
    .A(\memory[12][6] ),
    .B(_01575_),
    .Y(_02427_)
  );
  NAND _10586_ (
    .A(\memory[7][6] ),
    .B(_01517_),
    .Y(_02428_)
  );
  AND _10587_ (
    .A(_02427_),
    .B(_02428_),
    .Y(_02429_)
  );
  NAND _10588_ (
    .A(\memory[27][6] ),
    .B(_01484_),
    .Y(_02430_)
  );
  NAND _10589_ (
    .A(\memory[16][6] ),
    .B(_01501_),
    .Y(_02431_)
  );
  AND _10590_ (
    .A(_02430_),
    .B(_02431_),
    .Y(_02432_)
  );
  AND _10591_ (
    .A(_02429_),
    .B(_02432_),
    .Y(_02433_)
  );
  NAND _10592_ (
    .A(\memory[26][6] ),
    .B(_01559_),
    .Y(_02434_)
  );
  NAND _10593_ (
    .A(\memory[22][6] ),
    .B(_01474_),
    .Y(_02435_)
  );
  AND _10594_ (
    .A(_02434_),
    .B(_02435_),
    .Y(_02436_)
  );
  NAND _10595_ (
    .A(\memory[8][6] ),
    .B(_01538_),
    .Y(_02437_)
  );
  NAND _10596_ (
    .A(\memory[19][6] ),
    .B(_01582_),
    .Y(_02438_)
  );
  AND _10597_ (
    .A(_02437_),
    .B(_02438_),
    .Y(_02439_)
  );
  AND _10598_ (
    .A(_02436_),
    .B(_02439_),
    .Y(_02440_)
  );
  AND _10599_ (
    .A(_02433_),
    .B(_02440_),
    .Y(_02441_)
  );
  AND _10600_ (
    .A(_02426_),
    .B(_02441_),
    .Y(_02442_)
  );
  NAND _10601_ (
    .A(\memory[20][6] ),
    .B(_01534_),
    .Y(_02443_)
  );
  NAND _10602_ (
    .A(\memory[24][6] ),
    .B(_01546_),
    .Y(_02444_)
  );
  AND _10603_ (
    .A(_02443_),
    .B(_02444_),
    .Y(_02445_)
  );
  NAND _10604_ (
    .A(\memory[10][6] ),
    .B(_01495_),
    .Y(_02446_)
  );
  NAND _10605_ (
    .A(\memory[14][6] ),
    .B(_01520_),
    .Y(_02447_)
  );
  AND _10606_ (
    .A(_02446_),
    .B(_02447_),
    .Y(_02448_)
  );
  AND _10607_ (
    .A(_02445_),
    .B(_02448_),
    .Y(_02449_)
  );
  NAND _10608_ (
    .A(\memory[2][6] ),
    .B(_01570_),
    .Y(_02450_)
  );
  NAND _10609_ (
    .A(\memory[4][6] ),
    .B(_01513_),
    .Y(_02451_)
  );
  AND _10610_ (
    .A(_02450_),
    .B(_02451_),
    .Y(_02452_)
  );
  NAND _10611_ (
    .A(\memory[9][6] ),
    .B(_01527_),
    .Y(_02453_)
  );
  NAND _10612_ (
    .A(\memory[18][6] ),
    .B(_01479_),
    .Y(_02454_)
  );
  AND _10613_ (
    .A(_02453_),
    .B(_02454_),
    .Y(_02455_)
  );
  AND _10614_ (
    .A(_02452_),
    .B(_02455_),
    .Y(_02456_)
  );
  AND _10615_ (
    .A(_02449_),
    .B(_02456_),
    .Y(_02457_)
  );
  NAND _10616_ (
    .A(\memory[3][6] ),
    .B(_01453_),
    .Y(_02458_)
  );
  NAND _10617_ (
    .A(\memory[13][6] ),
    .B(_01458_),
    .Y(_02459_)
  );
  AND _10618_ (
    .A(_02458_),
    .B(_02459_),
    .Y(_02460_)
  );
  NAND _10619_ (
    .A(\memory[17][6] ),
    .B(_01567_),
    .Y(_02461_)
  );
  NAND _10620_ (
    .A(\memory[31][6] ),
    .B(_01491_),
    .Y(_02462_)
  );
  AND _10621_ (
    .A(_02461_),
    .B(_02462_),
    .Y(_02463_)
  );
  AND _10622_ (
    .A(_02460_),
    .B(_02463_),
    .Y(_02464_)
  );
  NAND _10623_ (
    .A(\memory[11][6] ),
    .B(_01578_),
    .Y(_02465_)
  );
  NAND _10624_ (
    .A(\memory[23][6] ),
    .B(_01469_),
    .Y(_02466_)
  );
  AND _10625_ (
    .A(_02465_),
    .B(_02466_),
    .Y(_02467_)
  );
  NAND _10626_ (
    .A(\memory[25][6] ),
    .B(_01550_),
    .Y(_02468_)
  );
  NAND _10627_ (
    .A(\memory[28][6] ),
    .B(_01563_),
    .Y(_02469_)
  );
  AND _10628_ (
    .A(_02468_),
    .B(_02469_),
    .Y(_02470_)
  );
  AND _10629_ (
    .A(_02467_),
    .B(_02470_),
    .Y(_02471_)
  );
  AND _10630_ (
    .A(_02464_),
    .B(_02471_),
    .Y(_02472_)
  );
  AND _10631_ (
    .A(_02457_),
    .B(_02472_),
    .Y(_02473_)
  );
  NAND _10632_ (
    .A(_02442_),
    .B(_02473_),
    .Y(_02474_)
  );
  AND _10633_ (
    .A(MemRead_i),
    .B(_02474_),
    .Y(\data_o[14] )
  );
  NAND _10634_ (
    .A(\memory[2][7] ),
    .B(_01570_),
    .Y(_02475_)
  );
  NAND _10635_ (
    .A(\memory[17][7] ),
    .B(_01567_),
    .Y(_02476_)
  );
  AND _10636_ (
    .A(_02475_),
    .B(_02476_),
    .Y(_02477_)
  );
  NAND _10637_ (
    .A(\memory[20][7] ),
    .B(_01534_),
    .Y(_02478_)
  );
  NAND _10638_ (
    .A(\memory[9][7] ),
    .B(_01527_),
    .Y(_02479_)
  );
  AND _10639_ (
    .A(_02478_),
    .B(_02479_),
    .Y(_02480_)
  );
  AND _10640_ (
    .A(_02477_),
    .B(_02480_),
    .Y(_02481_)
  );
  NAND _10641_ (
    .A(\memory[13][7] ),
    .B(_01458_),
    .Y(_02482_)
  );
  NAND _10642_ (
    .A(\memory[14][7] ),
    .B(_01520_),
    .Y(_02483_)
  );
  AND _10643_ (
    .A(_02482_),
    .B(_02483_),
    .Y(_02484_)
  );
  NAND _10644_ (
    .A(\memory[8][7] ),
    .B(_01538_),
    .Y(_02485_)
  );
  NAND _10645_ (
    .A(\memory[15][7] ),
    .B(_01543_),
    .Y(_02486_)
  );
  AND _10646_ (
    .A(_02485_),
    .B(_02486_),
    .Y(_02487_)
  );
  AND _10647_ (
    .A(_02484_),
    .B(_02487_),
    .Y(_02488_)
  );
  AND _10648_ (
    .A(_02481_),
    .B(_02488_),
    .Y(_02489_)
  );
  NAND _10649_ (
    .A(\memory[27][7] ),
    .B(_01484_),
    .Y(_02490_)
  );
  NAND _10650_ (
    .A(\memory[0][7] ),
    .B(_01504_),
    .Y(_02491_)
  );
  AND _10651_ (
    .A(_02490_),
    .B(_02491_),
    .Y(_02492_)
  );
  NAND _10652_ (
    .A(\memory[6][7] ),
    .B(_01585_),
    .Y(_02493_)
  );
  NAND _10653_ (
    .A(\memory[3][7] ),
    .B(_01453_),
    .Y(_02494_)
  );
  AND _10654_ (
    .A(_02493_),
    .B(_02494_),
    .Y(_02495_)
  );
  AND _10655_ (
    .A(_02492_),
    .B(_02495_),
    .Y(_02496_)
  );
  NAND _10656_ (
    .A(\memory[23][7] ),
    .B(_01469_),
    .Y(_02497_)
  );
  NAND _10657_ (
    .A(\memory[26][7] ),
    .B(_01559_),
    .Y(_02498_)
  );
  AND _10658_ (
    .A(_02497_),
    .B(_02498_),
    .Y(_02499_)
  );
  NAND _10659_ (
    .A(\memory[24][7] ),
    .B(_01546_),
    .Y(_02500_)
  );
  NAND _10660_ (
    .A(\memory[19][7] ),
    .B(_01582_),
    .Y(_02501_)
  );
  AND _10661_ (
    .A(_02500_),
    .B(_02501_),
    .Y(_02502_)
  );
  AND _10662_ (
    .A(_02499_),
    .B(_02502_),
    .Y(_02503_)
  );
  AND _10663_ (
    .A(_02496_),
    .B(_02503_),
    .Y(_02504_)
  );
  AND _10664_ (
    .A(_02489_),
    .B(_02504_),
    .Y(_02505_)
  );
  NAND _10665_ (
    .A(\memory[18][7] ),
    .B(_01479_),
    .Y(_02506_)
  );
  NAND _10666_ (
    .A(\memory[4][7] ),
    .B(_01513_),
    .Y(_02507_)
  );
  AND _10667_ (
    .A(_02506_),
    .B(_02507_),
    .Y(_02508_)
  );
  NAND _10668_ (
    .A(\memory[31][7] ),
    .B(_01491_),
    .Y(_02509_)
  );
  NAND _10669_ (
    .A(\memory[29][7] ),
    .B(_01462_),
    .Y(_02510_)
  );
  AND _10670_ (
    .A(_02509_),
    .B(_02510_),
    .Y(_02511_)
  );
  AND _10671_ (
    .A(_02508_),
    .B(_02511_),
    .Y(_02512_)
  );
  NAND _10672_ (
    .A(\memory[25][7] ),
    .B(_01550_),
    .Y(_02513_)
  );
  NAND _10673_ (
    .A(\memory[22][7] ),
    .B(_01474_),
    .Y(_02514_)
  );
  AND _10674_ (
    .A(_02513_),
    .B(_02514_),
    .Y(_02515_)
  );
  NAND _10675_ (
    .A(\memory[12][7] ),
    .B(_01575_),
    .Y(_02516_)
  );
  NAND _10676_ (
    .A(\memory[7][7] ),
    .B(_01517_),
    .Y(_02517_)
  );
  AND _10677_ (
    .A(_02516_),
    .B(_02517_),
    .Y(_02518_)
  );
  AND _10678_ (
    .A(_02515_),
    .B(_02518_),
    .Y(_02519_)
  );
  AND _10679_ (
    .A(_02512_),
    .B(_02519_),
    .Y(_02520_)
  );
  NAND _10680_ (
    .A(\memory[16][7] ),
    .B(_01501_),
    .Y(_02521_)
  );
  NAND _10681_ (
    .A(\memory[11][7] ),
    .B(_01578_),
    .Y(_02522_)
  );
  AND _10682_ (
    .A(_02521_),
    .B(_02522_),
    .Y(_02523_)
  );
  NAND _10683_ (
    .A(\memory[5][7] ),
    .B(_01530_),
    .Y(_02524_)
  );
  NAND _10684_ (
    .A(\memory[10][7] ),
    .B(_01495_),
    .Y(_02525_)
  );
  AND _10685_ (
    .A(_02524_),
    .B(_02525_),
    .Y(_02526_)
  );
  AND _10686_ (
    .A(_02523_),
    .B(_02526_),
    .Y(_02527_)
  );
  NAND _10687_ (
    .A(\memory[21][7] ),
    .B(_01553_),
    .Y(_02528_)
  );
  NAND _10688_ (
    .A(\memory[28][7] ),
    .B(_01563_),
    .Y(_02529_)
  );
  AND _10689_ (
    .A(_02528_),
    .B(_02529_),
    .Y(_02530_)
  );
  NAND _10690_ (
    .A(\memory[1][7] ),
    .B(_01449_),
    .Y(_02531_)
  );
  NAND _10691_ (
    .A(\memory[30][7] ),
    .B(_01510_),
    .Y(_02532_)
  );
  AND _10692_ (
    .A(_02531_),
    .B(_02532_),
    .Y(_02533_)
  );
  AND _10693_ (
    .A(_02530_),
    .B(_02533_),
    .Y(_02534_)
  );
  AND _10694_ (
    .A(_02527_),
    .B(_02534_),
    .Y(_02535_)
  );
  AND _10695_ (
    .A(_02520_),
    .B(_02535_),
    .Y(_02536_)
  );
  NAND _10696_ (
    .A(_02505_),
    .B(_02536_),
    .Y(_02537_)
  );
  AND _10697_ (
    .A(MemRead_i),
    .B(_02537_),
    .Y(\data_o[15] )
  );
  NAND _10698_ (
    .A(\memory[12][0] ),
    .B(_01578_),
    .Y(_02538_)
  );
  NAND _10699_ (
    .A(\memory[28][0] ),
    .B(_01484_),
    .Y(_02539_)
  );
  AND _10700_ (
    .A(_02538_),
    .B(_02539_),
    .Y(_02540_)
  );
  NAND _10701_ (
    .A(\memory[17][0] ),
    .B(_01501_),
    .Y(_02541_)
  );
  NAND _10702_ (
    .A(\memory[16][0] ),
    .B(_01543_),
    .Y(_02542_)
  );
  AND _10703_ (
    .A(_02541_),
    .B(_02542_),
    .Y(_02543_)
  );
  AND _10704_ (
    .A(_02540_),
    .B(_02543_),
    .Y(_02544_)
  );
  NAND _10705_ (
    .A(\memory[8][0] ),
    .B(_01517_),
    .Y(_02545_)
  );
  NAND _10706_ (
    .A(\memory[2][0] ),
    .B(_01449_),
    .Y(_02546_)
  );
  AND _10707_ (
    .A(_02545_),
    .B(_02546_),
    .Y(_02547_)
  );
  NAND _10708_ (
    .A(\memory[30][0] ),
    .B(_01462_),
    .Y(_02548_)
  );
  NAND _10709_ (
    .A(\memory[31][0] ),
    .B(_01510_),
    .Y(_02549_)
  );
  AND _10710_ (
    .A(_02548_),
    .B(_02549_),
    .Y(_02550_)
  );
  AND _10711_ (
    .A(_02547_),
    .B(_02550_),
    .Y(_02551_)
  );
  AND _10712_ (
    .A(_02544_),
    .B(_02551_),
    .Y(_02552_)
  );
  NAND _10713_ (
    .A(\memory[1][0] ),
    .B(_01504_),
    .Y(_02553_)
  );
  NAND _10714_ (
    .A(\memory[27][0] ),
    .B(_01559_),
    .Y(_02554_)
  );
  AND _10715_ (
    .A(_02553_),
    .B(_02554_),
    .Y(_02555_)
  );
  NAND _10716_ (
    .A(\memory[23][0] ),
    .B(_01474_),
    .Y(_02556_)
  );
  NAND _10717_ (
    .A(\memory[15][0] ),
    .B(_01520_),
    .Y(_02557_)
  );
  AND _10718_ (
    .A(_02556_),
    .B(_02557_),
    .Y(_02558_)
  );
  AND _10719_ (
    .A(_02555_),
    .B(_02558_),
    .Y(_02559_)
  );
  NAND _10720_ (
    .A(\memory[21][0] ),
    .B(_01534_),
    .Y(_02560_)
  );
  NAND _10721_ (
    .A(\memory[24][0] ),
    .B(_01469_),
    .Y(_02561_)
  );
  AND _10722_ (
    .A(_02560_),
    .B(_02561_),
    .Y(_02562_)
  );
  NAND _10723_ (
    .A(\memory[18][0] ),
    .B(_01567_),
    .Y(_02563_)
  );
  NAND _10724_ (
    .A(\memory[11][0] ),
    .B(_01495_),
    .Y(_02564_)
  );
  AND _10725_ (
    .A(_02563_),
    .B(_02564_),
    .Y(_02565_)
  );
  AND _10726_ (
    .A(_02562_),
    .B(_02565_),
    .Y(_02566_)
  );
  AND _10727_ (
    .A(_02559_),
    .B(_02566_),
    .Y(_02567_)
  );
  AND _10728_ (
    .A(_02552_),
    .B(_02567_),
    .Y(_02568_)
  );
  NAND _10729_ (
    .A(\memory[25][0] ),
    .B(_01546_),
    .Y(_02569_)
  );
  NAND _10730_ (
    .A(\memory[22][0] ),
    .B(_01553_),
    .Y(_02570_)
  );
  AND _10731_ (
    .A(_02569_),
    .B(_02570_),
    .Y(_02571_)
  );
  NAND _10732_ (
    .A(\memory[14][0] ),
    .B(_01458_),
    .Y(_02572_)
  );
  NAND _10733_ (
    .A(\memory[29][0] ),
    .B(_01563_),
    .Y(_02573_)
  );
  AND _10734_ (
    .A(_02572_),
    .B(_02573_),
    .Y(_02574_)
  );
  AND _10735_ (
    .A(_02571_),
    .B(_02574_),
    .Y(_02575_)
  );
  NAND _10736_ (
    .A(\memory[19][0] ),
    .B(_01479_),
    .Y(_02576_)
  );
  NAND _10737_ (
    .A(\memory[7][0] ),
    .B(_01585_),
    .Y(_02577_)
  );
  AND _10738_ (
    .A(_02576_),
    .B(_02577_),
    .Y(_02578_)
  );
  NAND _10739_ (
    .A(\memory[3][0] ),
    .B(_01570_),
    .Y(_02579_)
  );
  NAND _10740_ (
    .A(\memory[13][0] ),
    .B(_01575_),
    .Y(_02580_)
  );
  AND _10741_ (
    .A(_02579_),
    .B(_02580_),
    .Y(_02581_)
  );
  AND _10742_ (
    .A(_02578_),
    .B(_02581_),
    .Y(_02582_)
  );
  AND _10743_ (
    .A(_02575_),
    .B(_02582_),
    .Y(_02583_)
  );
  NAND _10744_ (
    .A(\memory[26][0] ),
    .B(_01550_),
    .Y(_02584_)
  );
  NAND _10745_ (
    .A(\memory[0][0] ),
    .B(_01491_),
    .Y(_02585_)
  );
  AND _10746_ (
    .A(_02584_),
    .B(_02585_),
    .Y(_02586_)
  );
  NAND _10747_ (
    .A(\memory[20][0] ),
    .B(_01582_),
    .Y(_02587_)
  );
  NAND _10748_ (
    .A(\memory[9][0] ),
    .B(_01538_),
    .Y(_02588_)
  );
  AND _10749_ (
    .A(_02587_),
    .B(_02588_),
    .Y(_02589_)
  );
  AND _10750_ (
    .A(_02586_),
    .B(_02589_),
    .Y(_02590_)
  );
  NAND _10751_ (
    .A(\memory[5][0] ),
    .B(_01513_),
    .Y(_02591_)
  );
  NAND _10752_ (
    .A(\memory[6][0] ),
    .B(_01530_),
    .Y(_02592_)
  );
  AND _10753_ (
    .A(_02591_),
    .B(_02592_),
    .Y(_02593_)
  );
  NAND _10754_ (
    .A(\memory[4][0] ),
    .B(_01453_),
    .Y(_02594_)
  );
  NAND _10755_ (
    .A(\memory[10][0] ),
    .B(_01527_),
    .Y(_02595_)
  );
  AND _10756_ (
    .A(_02594_),
    .B(_02595_),
    .Y(_02596_)
  );
  AND _10757_ (
    .A(_02593_),
    .B(_02596_),
    .Y(_02597_)
  );
  AND _10758_ (
    .A(_02590_),
    .B(_02597_),
    .Y(_02598_)
  );
  AND _10759_ (
    .A(_02583_),
    .B(_02598_),
    .Y(_02599_)
  );
  NAND _10760_ (
    .A(_02568_),
    .B(_02599_),
    .Y(_02600_)
  );
  AND _10761_ (
    .A(MemRead_i),
    .B(_02600_),
    .Y(\data_o[16] )
  );
  NAND _10762_ (
    .A(\memory[19][1] ),
    .B(_01479_),
    .Y(_02601_)
  );
  NAND _10763_ (
    .A(\memory[28][1] ),
    .B(_01484_),
    .Y(_02602_)
  );
  AND _10764_ (
    .A(_02601_),
    .B(_02602_),
    .Y(_02603_)
  );
  NAND _10765_ (
    .A(\memory[23][1] ),
    .B(_01474_),
    .Y(_02604_)
  );
  NAND _10766_ (
    .A(\memory[6][1] ),
    .B(_01530_),
    .Y(_02605_)
  );
  AND _10767_ (
    .A(_02604_),
    .B(_02605_),
    .Y(_02606_)
  );
  AND _10768_ (
    .A(_02603_),
    .B(_02606_),
    .Y(_02607_)
  );
  NAND _10769_ (
    .A(\memory[15][1] ),
    .B(_01520_),
    .Y(_02608_)
  );
  NAND _10770_ (
    .A(\memory[2][1] ),
    .B(_01449_),
    .Y(_02609_)
  );
  AND _10771_ (
    .A(_02608_),
    .B(_02609_),
    .Y(_02610_)
  );
  NAND _10772_ (
    .A(\memory[14][1] ),
    .B(_01458_),
    .Y(_02611_)
  );
  NAND _10773_ (
    .A(\memory[29][1] ),
    .B(_01563_),
    .Y(_02612_)
  );
  AND _10774_ (
    .A(_02611_),
    .B(_02612_),
    .Y(_02613_)
  );
  AND _10775_ (
    .A(_02610_),
    .B(_02613_),
    .Y(_02614_)
  );
  AND _10776_ (
    .A(_02607_),
    .B(_02614_),
    .Y(_02615_)
  );
  NAND _10777_ (
    .A(\memory[8][1] ),
    .B(_01517_),
    .Y(_02616_)
  );
  NAND _10778_ (
    .A(\memory[27][1] ),
    .B(_01559_),
    .Y(_02617_)
  );
  AND _10779_ (
    .A(_02616_),
    .B(_02617_),
    .Y(_02618_)
  );
  NAND _10780_ (
    .A(\memory[11][1] ),
    .B(_01495_),
    .Y(_02619_)
  );
  NAND _10781_ (
    .A(\memory[16][1] ),
    .B(_01543_),
    .Y(_02620_)
  );
  AND _10782_ (
    .A(_02619_),
    .B(_02620_),
    .Y(_02621_)
  );
  AND _10783_ (
    .A(_02618_),
    .B(_02621_),
    .Y(_02622_)
  );
  NAND _10784_ (
    .A(\memory[9][1] ),
    .B(_01538_),
    .Y(_02623_)
  );
  NAND _10785_ (
    .A(\memory[7][1] ),
    .B(_01585_),
    .Y(_02624_)
  );
  AND _10786_ (
    .A(_02623_),
    .B(_02624_),
    .Y(_02625_)
  );
  NAND _10787_ (
    .A(\memory[20][1] ),
    .B(_01582_),
    .Y(_02626_)
  );
  NAND _10788_ (
    .A(\memory[10][1] ),
    .B(_01527_),
    .Y(_02627_)
  );
  AND _10789_ (
    .A(_02626_),
    .B(_02627_),
    .Y(_02628_)
  );
  AND _10790_ (
    .A(_02625_),
    .B(_02628_),
    .Y(_02629_)
  );
  AND _10791_ (
    .A(_02622_),
    .B(_02629_),
    .Y(_02630_)
  );
  AND _10792_ (
    .A(_02615_),
    .B(_02630_),
    .Y(_02631_)
  );
  NAND _10793_ (
    .A(\memory[5][1] ),
    .B(_01513_),
    .Y(_02632_)
  );
  NAND _10794_ (
    .A(\memory[1][1] ),
    .B(_01504_),
    .Y(_02633_)
  );
  AND _10795_ (
    .A(_02632_),
    .B(_02633_),
    .Y(_02634_)
  );
  NAND _10796_ (
    .A(\memory[30][1] ),
    .B(_01462_),
    .Y(_02635_)
  );
  NAND _10797_ (
    .A(\memory[31][1] ),
    .B(_01510_),
    .Y(_02636_)
  );
  AND _10798_ (
    .A(_02635_),
    .B(_02636_),
    .Y(_02637_)
  );
  AND _10799_ (
    .A(_02634_),
    .B(_02637_),
    .Y(_02638_)
  );
  NAND _10800_ (
    .A(\memory[24][1] ),
    .B(_01469_),
    .Y(_02639_)
  );
  NAND _10801_ (
    .A(\memory[18][1] ),
    .B(_01567_),
    .Y(_02640_)
  );
  AND _10802_ (
    .A(_02639_),
    .B(_02640_),
    .Y(_02641_)
  );
  NAND _10803_ (
    .A(\memory[22][1] ),
    .B(_01553_),
    .Y(_02642_)
  );
  NAND _10804_ (
    .A(\memory[13][1] ),
    .B(_01575_),
    .Y(_02643_)
  );
  AND _10805_ (
    .A(_02642_),
    .B(_02643_),
    .Y(_02644_)
  );
  AND _10806_ (
    .A(_02641_),
    .B(_02644_),
    .Y(_02645_)
  );
  AND _10807_ (
    .A(_02638_),
    .B(_02645_),
    .Y(_02646_)
  );
  NAND _10808_ (
    .A(\memory[26][1] ),
    .B(_01550_),
    .Y(_02647_)
  );
  NAND _10809_ (
    .A(\memory[0][1] ),
    .B(_01491_),
    .Y(_02648_)
  );
  AND _10810_ (
    .A(_02647_),
    .B(_02648_),
    .Y(_02649_)
  );
  NAND _10811_ (
    .A(\memory[12][1] ),
    .B(_01578_),
    .Y(_02650_)
  );
  NAND _10812_ (
    .A(\memory[21][1] ),
    .B(_01534_),
    .Y(_02651_)
  );
  AND _10813_ (
    .A(_02650_),
    .B(_02651_),
    .Y(_02652_)
  );
  AND _10814_ (
    .A(_02649_),
    .B(_02652_),
    .Y(_02653_)
  );
  NAND _10815_ (
    .A(\memory[3][1] ),
    .B(_01570_),
    .Y(_02654_)
  );
  NAND _10816_ (
    .A(\memory[4][1] ),
    .B(_01453_),
    .Y(_02655_)
  );
  AND _10817_ (
    .A(_02654_),
    .B(_02655_),
    .Y(_02656_)
  );
  NAND _10818_ (
    .A(\memory[17][1] ),
    .B(_01501_),
    .Y(_02657_)
  );
  NAND _10819_ (
    .A(\memory[25][1] ),
    .B(_01546_),
    .Y(_02658_)
  );
  AND _10820_ (
    .A(_02657_),
    .B(_02658_),
    .Y(_02659_)
  );
  AND _10821_ (
    .A(_02656_),
    .B(_02659_),
    .Y(_02660_)
  );
  AND _10822_ (
    .A(_02653_),
    .B(_02660_),
    .Y(_02661_)
  );
  AND _10823_ (
    .A(_02646_),
    .B(_02661_),
    .Y(_02662_)
  );
  NAND _10824_ (
    .A(_02631_),
    .B(_02662_),
    .Y(_02663_)
  );
  AND _10825_ (
    .A(MemRead_i),
    .B(_02663_),
    .Y(\data_o[17] )
  );
  NAND _10826_ (
    .A(\memory[0][2] ),
    .B(_01491_),
    .Y(_02664_)
  );
  NAND _10827_ (
    .A(\memory[30][2] ),
    .B(_01462_),
    .Y(_02665_)
  );
  AND _10828_ (
    .A(_02664_),
    .B(_02665_),
    .Y(_02666_)
  );
  NAND _10829_ (
    .A(\memory[26][2] ),
    .B(_01550_),
    .Y(_02667_)
  );
  NAND _10830_ (
    .A(\memory[27][2] ),
    .B(_01559_),
    .Y(_02668_)
  );
  AND _10831_ (
    .A(_02667_),
    .B(_02668_),
    .Y(_02669_)
  );
  AND _10832_ (
    .A(_02666_),
    .B(_02669_),
    .Y(_02670_)
  );
  NAND _10833_ (
    .A(\memory[29][2] ),
    .B(_01563_),
    .Y(_02671_)
  );
  NAND _10834_ (
    .A(\memory[28][2] ),
    .B(_01484_),
    .Y(_02672_)
  );
  AND _10835_ (
    .A(_02671_),
    .B(_02672_),
    .Y(_02673_)
  );
  NAND _10836_ (
    .A(\memory[14][2] ),
    .B(_01458_),
    .Y(_02674_)
  );
  NAND _10837_ (
    .A(\memory[11][2] ),
    .B(_01495_),
    .Y(_02675_)
  );
  AND _10838_ (
    .A(_02674_),
    .B(_02675_),
    .Y(_02676_)
  );
  AND _10839_ (
    .A(_02673_),
    .B(_02676_),
    .Y(_02677_)
  );
  AND _10840_ (
    .A(_02670_),
    .B(_02677_),
    .Y(_02678_)
  );
  NAND _10841_ (
    .A(\memory[12][2] ),
    .B(_01578_),
    .Y(_02679_)
  );
  NAND _10842_ (
    .A(\memory[15][2] ),
    .B(_01520_),
    .Y(_02680_)
  );
  AND _10843_ (
    .A(_02679_),
    .B(_02680_),
    .Y(_02681_)
  );
  NAND _10844_ (
    .A(\memory[24][2] ),
    .B(_01469_),
    .Y(_02682_)
  );
  NAND _10845_ (
    .A(\memory[25][2] ),
    .B(_01546_),
    .Y(_02683_)
  );
  AND _10846_ (
    .A(_02682_),
    .B(_02683_),
    .Y(_02684_)
  );
  AND _10847_ (
    .A(_02681_),
    .B(_02684_),
    .Y(_02685_)
  );
  NAND _10848_ (
    .A(\memory[20][2] ),
    .B(_01582_),
    .Y(_02686_)
  );
  NAND _10849_ (
    .A(\memory[10][2] ),
    .B(_01527_),
    .Y(_02687_)
  );
  AND _10850_ (
    .A(_02686_),
    .B(_02687_),
    .Y(_02688_)
  );
  NAND _10851_ (
    .A(\memory[9][2] ),
    .B(_01538_),
    .Y(_02689_)
  );
  NAND _10852_ (
    .A(\memory[7][2] ),
    .B(_01585_),
    .Y(_02690_)
  );
  AND _10853_ (
    .A(_02689_),
    .B(_02690_),
    .Y(_02691_)
  );
  AND _10854_ (
    .A(_02688_),
    .B(_02691_),
    .Y(_02692_)
  );
  AND _10855_ (
    .A(_02685_),
    .B(_02692_),
    .Y(_02693_)
  );
  AND _10856_ (
    .A(_02678_),
    .B(_02693_),
    .Y(_02694_)
  );
  NAND _10857_ (
    .A(\memory[5][2] ),
    .B(_01513_),
    .Y(_02695_)
  );
  NAND _10858_ (
    .A(\memory[4][2] ),
    .B(_01453_),
    .Y(_02696_)
  );
  AND _10859_ (
    .A(_02695_),
    .B(_02696_),
    .Y(_02697_)
  );
  NAND _10860_ (
    .A(\memory[16][2] ),
    .B(_01543_),
    .Y(_02698_)
  );
  NAND _10861_ (
    .A(\memory[17][2] ),
    .B(_01501_),
    .Y(_02699_)
  );
  AND _10862_ (
    .A(_02698_),
    .B(_02699_),
    .Y(_02700_)
  );
  AND _10863_ (
    .A(_02697_),
    .B(_02700_),
    .Y(_02701_)
  );
  NAND _10864_ (
    .A(\memory[3][2] ),
    .B(_01570_),
    .Y(_02702_)
  );
  NAND _10865_ (
    .A(\memory[1][2] ),
    .B(_01504_),
    .Y(_02703_)
  );
  AND _10866_ (
    .A(_02702_),
    .B(_02703_),
    .Y(_02704_)
  );
  NAND _10867_ (
    .A(\memory[13][2] ),
    .B(_01575_),
    .Y(_02705_)
  );
  NAND _10868_ (
    .A(\memory[6][2] ),
    .B(_01530_),
    .Y(_02706_)
  );
  AND _10869_ (
    .A(_02705_),
    .B(_02706_),
    .Y(_02707_)
  );
  AND _10870_ (
    .A(_02704_),
    .B(_02707_),
    .Y(_02708_)
  );
  AND _10871_ (
    .A(_02701_),
    .B(_02708_),
    .Y(_02709_)
  );
  NAND _10872_ (
    .A(\memory[31][2] ),
    .B(_01510_),
    .Y(_02710_)
  );
  NAND _10873_ (
    .A(\memory[2][2] ),
    .B(_01449_),
    .Y(_02711_)
  );
  AND _10874_ (
    .A(_02710_),
    .B(_02711_),
    .Y(_02712_)
  );
  NAND _10875_ (
    .A(\memory[19][2] ),
    .B(_01479_),
    .Y(_02713_)
  );
  NAND _10876_ (
    .A(\memory[22][2] ),
    .B(_01553_),
    .Y(_02714_)
  );
  AND _10877_ (
    .A(_02713_),
    .B(_02714_),
    .Y(_02715_)
  );
  AND _10878_ (
    .A(_02712_),
    .B(_02715_),
    .Y(_02716_)
  );
  NAND _10879_ (
    .A(\memory[8][2] ),
    .B(_01517_),
    .Y(_02717_)
  );
  NAND _10880_ (
    .A(\memory[23][2] ),
    .B(_01474_),
    .Y(_02718_)
  );
  AND _10881_ (
    .A(_02717_),
    .B(_02718_),
    .Y(_02719_)
  );
  NAND _10882_ (
    .A(\memory[18][2] ),
    .B(_01567_),
    .Y(_02720_)
  );
  NAND _10883_ (
    .A(\memory[21][2] ),
    .B(_01534_),
    .Y(_02721_)
  );
  AND _10884_ (
    .A(_02720_),
    .B(_02721_),
    .Y(_02722_)
  );
  AND _10885_ (
    .A(_02719_),
    .B(_02722_),
    .Y(_02723_)
  );
  AND _10886_ (
    .A(_02716_),
    .B(_02723_),
    .Y(_02724_)
  );
  AND _10887_ (
    .A(_02709_),
    .B(_02724_),
    .Y(_02725_)
  );
  NAND _10888_ (
    .A(_02694_),
    .B(_02725_),
    .Y(_02726_)
  );
  AND _10889_ (
    .A(MemRead_i),
    .B(_02726_),
    .Y(\data_o[18] )
  );
  NAND _10890_ (
    .A(\memory[5][3] ),
    .B(_01513_),
    .Y(_02727_)
  );
  NAND _10891_ (
    .A(\memory[1][3] ),
    .B(_01504_),
    .Y(_02728_)
  );
  AND _10892_ (
    .A(_02727_),
    .B(_02728_),
    .Y(_02729_)
  );
  NAND _10893_ (
    .A(\memory[22][3] ),
    .B(_01553_),
    .Y(_02730_)
  );
  NAND _10894_ (
    .A(\memory[10][3] ),
    .B(_01527_),
    .Y(_02731_)
  );
  AND _10895_ (
    .A(_02730_),
    .B(_02731_),
    .Y(_02732_)
  );
  AND _10896_ (
    .A(_02729_),
    .B(_02732_),
    .Y(_02733_)
  );
  NAND _10897_ (
    .A(\memory[21][3] ),
    .B(_01534_),
    .Y(_02734_)
  );
  NAND _10898_ (
    .A(\memory[23][3] ),
    .B(_01474_),
    .Y(_02735_)
  );
  AND _10899_ (
    .A(_02734_),
    .B(_02735_),
    .Y(_02736_)
  );
  NAND _10900_ (
    .A(\memory[6][3] ),
    .B(_01530_),
    .Y(_02737_)
  );
  NAND _10901_ (
    .A(\memory[7][3] ),
    .B(_01585_),
    .Y(_02738_)
  );
  AND _10902_ (
    .A(_02737_),
    .B(_02738_),
    .Y(_02739_)
  );
  AND _10903_ (
    .A(_02736_),
    .B(_02739_),
    .Y(_02740_)
  );
  AND _10904_ (
    .A(_02733_),
    .B(_02740_),
    .Y(_02741_)
  );
  NAND _10905_ (
    .A(\memory[3][3] ),
    .B(_01570_),
    .Y(_02742_)
  );
  NAND _10906_ (
    .A(\memory[9][3] ),
    .B(_01538_),
    .Y(_02743_)
  );
  AND _10907_ (
    .A(_02742_),
    .B(_02743_),
    .Y(_02744_)
  );
  NAND _10908_ (
    .A(\memory[24][3] ),
    .B(_01469_),
    .Y(_02745_)
  );
  NAND _10909_ (
    .A(\memory[11][3] ),
    .B(_01495_),
    .Y(_02746_)
  );
  AND _10910_ (
    .A(_02745_),
    .B(_02746_),
    .Y(_02747_)
  );
  AND _10911_ (
    .A(_02744_),
    .B(_02747_),
    .Y(_02748_)
  );
  NAND _10912_ (
    .A(\memory[27][3] ),
    .B(_01559_),
    .Y(_02749_)
  );
  NAND _10913_ (
    .A(\memory[26][3] ),
    .B(_01550_),
    .Y(_02750_)
  );
  AND _10914_ (
    .A(_02749_),
    .B(_02750_),
    .Y(_02751_)
  );
  NAND _10915_ (
    .A(\memory[18][3] ),
    .B(_01567_),
    .Y(_02752_)
  );
  NAND _10916_ (
    .A(\memory[4][3] ),
    .B(_01453_),
    .Y(_02753_)
  );
  AND _10917_ (
    .A(_02752_),
    .B(_02753_),
    .Y(_02754_)
  );
  AND _10918_ (
    .A(_02751_),
    .B(_02754_),
    .Y(_02755_)
  );
  AND _10919_ (
    .A(_02748_),
    .B(_02755_),
    .Y(_02756_)
  );
  AND _10920_ (
    .A(_02741_),
    .B(_02756_),
    .Y(_02757_)
  );
  NAND _10921_ (
    .A(\memory[0][3] ),
    .B(_01491_),
    .Y(_02758_)
  );
  NAND _10922_ (
    .A(\memory[15][3] ),
    .B(_01520_),
    .Y(_02759_)
  );
  AND _10923_ (
    .A(_02758_),
    .B(_02759_),
    .Y(_02760_)
  );
  NAND _10924_ (
    .A(\memory[17][3] ),
    .B(_01501_),
    .Y(_02761_)
  );
  NAND _10925_ (
    .A(\memory[29][3] ),
    .B(_01563_),
    .Y(_02762_)
  );
  AND _10926_ (
    .A(_02761_),
    .B(_02762_),
    .Y(_02763_)
  );
  AND _10927_ (
    .A(_02760_),
    .B(_02763_),
    .Y(_02764_)
  );
  NAND _10928_ (
    .A(\memory[28][3] ),
    .B(_01484_),
    .Y(_02765_)
  );
  NAND _10929_ (
    .A(\memory[30][3] ),
    .B(_01462_),
    .Y(_02766_)
  );
  AND _10930_ (
    .A(_02765_),
    .B(_02766_),
    .Y(_02767_)
  );
  NAND _10931_ (
    .A(\memory[13][3] ),
    .B(_01575_),
    .Y(_02768_)
  );
  NAND _10932_ (
    .A(\memory[14][3] ),
    .B(_01458_),
    .Y(_02769_)
  );
  AND _10933_ (
    .A(_02768_),
    .B(_02769_),
    .Y(_02770_)
  );
  AND _10934_ (
    .A(_02767_),
    .B(_02770_),
    .Y(_02771_)
  );
  AND _10935_ (
    .A(_02764_),
    .B(_02771_),
    .Y(_02772_)
  );
  NAND _10936_ (
    .A(\memory[12][3] ),
    .B(_01578_),
    .Y(_02773_)
  );
  NAND _10937_ (
    .A(\memory[2][3] ),
    .B(_01449_),
    .Y(_02774_)
  );
  AND _10938_ (
    .A(_02773_),
    .B(_02774_),
    .Y(_02775_)
  );
  NAND _10939_ (
    .A(\memory[19][3] ),
    .B(_01479_),
    .Y(_02776_)
  );
  NAND _10940_ (
    .A(\memory[8][3] ),
    .B(_01517_),
    .Y(_02777_)
  );
  AND _10941_ (
    .A(_02776_),
    .B(_02777_),
    .Y(_02778_)
  );
  AND _10942_ (
    .A(_02775_),
    .B(_02778_),
    .Y(_02779_)
  );
  NAND _10943_ (
    .A(\memory[16][3] ),
    .B(_01543_),
    .Y(_02780_)
  );
  NAND _10944_ (
    .A(\memory[25][3] ),
    .B(_01546_),
    .Y(_02781_)
  );
  AND _10945_ (
    .A(_02780_),
    .B(_02781_),
    .Y(_02782_)
  );
  NAND _10946_ (
    .A(\memory[20][3] ),
    .B(_01582_),
    .Y(_02783_)
  );
  NAND _10947_ (
    .A(\memory[31][3] ),
    .B(_01510_),
    .Y(_02784_)
  );
  AND _10948_ (
    .A(_02783_),
    .B(_02784_),
    .Y(_02785_)
  );
  AND _10949_ (
    .A(_02782_),
    .B(_02785_),
    .Y(_02786_)
  );
  AND _10950_ (
    .A(_02779_),
    .B(_02786_),
    .Y(_02787_)
  );
  AND _10951_ (
    .A(_02772_),
    .B(_02787_),
    .Y(_02788_)
  );
  NAND _10952_ (
    .A(_02757_),
    .B(_02788_),
    .Y(_02789_)
  );
  AND _10953_ (
    .A(MemRead_i),
    .B(_02789_),
    .Y(\data_o[19] )
  );
  NAND _10954_ (
    .A(\memory[10][4] ),
    .B(_01527_),
    .Y(_02790_)
  );
  NAND _10955_ (
    .A(\memory[26][4] ),
    .B(_01550_),
    .Y(_02791_)
  );
  AND _10956_ (
    .A(_02790_),
    .B(_02791_),
    .Y(_02792_)
  );
  NAND _10957_ (
    .A(\memory[30][4] ),
    .B(_01462_),
    .Y(_02793_)
  );
  NAND _10958_ (
    .A(\memory[0][4] ),
    .B(_01491_),
    .Y(_02794_)
  );
  AND _10959_ (
    .A(_02793_),
    .B(_02794_),
    .Y(_02795_)
  );
  AND _10960_ (
    .A(_02792_),
    .B(_02795_),
    .Y(_02796_)
  );
  NAND _10961_ (
    .A(\memory[15][4] ),
    .B(_01520_),
    .Y(_02797_)
  );
  NAND _10962_ (
    .A(\memory[14][4] ),
    .B(_01458_),
    .Y(_02798_)
  );
  AND _10963_ (
    .A(_02797_),
    .B(_02798_),
    .Y(_02799_)
  );
  NAND _10964_ (
    .A(\memory[23][4] ),
    .B(_01474_),
    .Y(_02800_)
  );
  NAND _10965_ (
    .A(\memory[8][4] ),
    .B(_01517_),
    .Y(_02801_)
  );
  AND _10966_ (
    .A(_02800_),
    .B(_02801_),
    .Y(_02802_)
  );
  AND _10967_ (
    .A(_02799_),
    .B(_02802_),
    .Y(_02803_)
  );
  AND _10968_ (
    .A(_02796_),
    .B(_02803_),
    .Y(_02804_)
  );
  NAND _10969_ (
    .A(\memory[3][4] ),
    .B(_01570_),
    .Y(_02805_)
  );
  NAND _10970_ (
    .A(\memory[13][4] ),
    .B(_01575_),
    .Y(_02806_)
  );
  AND _10971_ (
    .A(_02805_),
    .B(_02806_),
    .Y(_02807_)
  );
  NAND _10972_ (
    .A(\memory[1][4] ),
    .B(_01504_),
    .Y(_02808_)
  );
  NAND _10973_ (
    .A(\memory[4][4] ),
    .B(_01453_),
    .Y(_02809_)
  );
  AND _10974_ (
    .A(_02808_),
    .B(_02809_),
    .Y(_02810_)
  );
  AND _10975_ (
    .A(_02807_),
    .B(_02810_),
    .Y(_02811_)
  );
  NAND _10976_ (
    .A(\memory[27][4] ),
    .B(_01559_),
    .Y(_02812_)
  );
  NAND _10977_ (
    .A(\memory[31][4] ),
    .B(_01510_),
    .Y(_02813_)
  );
  AND _10978_ (
    .A(_02812_),
    .B(_02813_),
    .Y(_02814_)
  );
  NAND _10979_ (
    .A(\memory[24][4] ),
    .B(_01469_),
    .Y(_02815_)
  );
  NAND _10980_ (
    .A(\memory[29][4] ),
    .B(_01563_),
    .Y(_02816_)
  );
  AND _10981_ (
    .A(_02815_),
    .B(_02816_),
    .Y(_02817_)
  );
  AND _10982_ (
    .A(_02814_),
    .B(_02817_),
    .Y(_02818_)
  );
  AND _10983_ (
    .A(_02811_),
    .B(_02818_),
    .Y(_02819_)
  );
  AND _10984_ (
    .A(_02804_),
    .B(_02819_),
    .Y(_02820_)
  );
  NAND _10985_ (
    .A(\memory[5][4] ),
    .B(_01513_),
    .Y(_02821_)
  );
  NAND _10986_ (
    .A(\memory[6][4] ),
    .B(_01530_),
    .Y(_02822_)
  );
  AND _10987_ (
    .A(_02821_),
    .B(_02822_),
    .Y(_02823_)
  );
  NAND _10988_ (
    .A(\memory[28][4] ),
    .B(_01484_),
    .Y(_02824_)
  );
  NAND _10989_ (
    .A(\memory[2][4] ),
    .B(_01449_),
    .Y(_02825_)
  );
  AND _10990_ (
    .A(_02824_),
    .B(_02825_),
    .Y(_02826_)
  );
  AND _10991_ (
    .A(_02823_),
    .B(_02826_),
    .Y(_02827_)
  );
  NAND _10992_ (
    .A(\memory[21][4] ),
    .B(_01534_),
    .Y(_02828_)
  );
  NAND _10993_ (
    .A(\memory[20][4] ),
    .B(_01582_),
    .Y(_02829_)
  );
  AND _10994_ (
    .A(_02828_),
    .B(_02829_),
    .Y(_02830_)
  );
  NAND _10995_ (
    .A(\memory[17][4] ),
    .B(_01501_),
    .Y(_02831_)
  );
  NAND _10996_ (
    .A(\memory[12][4] ),
    .B(_01578_),
    .Y(_02832_)
  );
  AND _10997_ (
    .A(_02831_),
    .B(_02832_),
    .Y(_02833_)
  );
  AND _10998_ (
    .A(_02830_),
    .B(_02833_),
    .Y(_02834_)
  );
  AND _10999_ (
    .A(_02827_),
    .B(_02834_),
    .Y(_02835_)
  );
  NAND _11000_ (
    .A(\memory[19][4] ),
    .B(_01479_),
    .Y(_02836_)
  );
  NAND _11001_ (
    .A(\memory[7][4] ),
    .B(_01585_),
    .Y(_02837_)
  );
  AND _11002_ (
    .A(_02836_),
    .B(_02837_),
    .Y(_02838_)
  );
  NAND _11003_ (
    .A(\memory[9][4] ),
    .B(_01538_),
    .Y(_02839_)
  );
  NAND _11004_ (
    .A(\memory[16][4] ),
    .B(_01543_),
    .Y(_02840_)
  );
  AND _11005_ (
    .A(_02839_),
    .B(_02840_),
    .Y(_02841_)
  );
  AND _11006_ (
    .A(_02838_),
    .B(_02841_),
    .Y(_02842_)
  );
  NAND _11007_ (
    .A(\memory[25][4] ),
    .B(_01546_),
    .Y(_02843_)
  );
  NAND _11008_ (
    .A(\memory[22][4] ),
    .B(_01553_),
    .Y(_02844_)
  );
  AND _11009_ (
    .A(_02843_),
    .B(_02844_),
    .Y(_02845_)
  );
  NAND _11010_ (
    .A(\memory[11][4] ),
    .B(_01495_),
    .Y(_02846_)
  );
  NAND _11011_ (
    .A(\memory[18][4] ),
    .B(_01567_),
    .Y(_02847_)
  );
  AND _11012_ (
    .A(_02846_),
    .B(_02847_),
    .Y(_02848_)
  );
  AND _11013_ (
    .A(_02845_),
    .B(_02848_),
    .Y(_02849_)
  );
  AND _11014_ (
    .A(_02842_),
    .B(_02849_),
    .Y(_02850_)
  );
  AND _11015_ (
    .A(_02835_),
    .B(_02850_),
    .Y(_02851_)
  );
  NAND _11016_ (
    .A(_02820_),
    .B(_02851_),
    .Y(_02852_)
  );
  AND _11017_ (
    .A(MemRead_i),
    .B(_02852_),
    .Y(\data_o[20] )
  );
  NAND _11018_ (
    .A(\memory[8][5] ),
    .B(_01517_),
    .Y(_02853_)
  );
  NAND _11019_ (
    .A(\memory[18][5] ),
    .B(_01567_),
    .Y(_02854_)
  );
  AND _11020_ (
    .A(_02853_),
    .B(_02854_),
    .Y(_02855_)
  );
  NAND _11021_ (
    .A(\memory[20][5] ),
    .B(_01582_),
    .Y(_02856_)
  );
  NAND _11022_ (
    .A(\memory[31][5] ),
    .B(_01510_),
    .Y(_02857_)
  );
  AND _11023_ (
    .A(_02856_),
    .B(_02857_),
    .Y(_02858_)
  );
  AND _11024_ (
    .A(_02855_),
    .B(_02858_),
    .Y(_02859_)
  );
  NAND _11025_ (
    .A(\memory[5][5] ),
    .B(_01513_),
    .Y(_02860_)
  );
  NAND _11026_ (
    .A(\memory[10][5] ),
    .B(_01527_),
    .Y(_02861_)
  );
  AND _11027_ (
    .A(_02860_),
    .B(_02861_),
    .Y(_02862_)
  );
  NAND _11028_ (
    .A(\memory[13][5] ),
    .B(_01575_),
    .Y(_02863_)
  );
  NAND _11029_ (
    .A(\memory[27][5] ),
    .B(_01559_),
    .Y(_02864_)
  );
  AND _11030_ (
    .A(_02863_),
    .B(_02864_),
    .Y(_02865_)
  );
  AND _11031_ (
    .A(_02862_),
    .B(_02865_),
    .Y(_02866_)
  );
  AND _11032_ (
    .A(_02859_),
    .B(_02866_),
    .Y(_02867_)
  );
  NAND _11033_ (
    .A(\memory[1][5] ),
    .B(_01504_),
    .Y(_02868_)
  );
  NAND _11034_ (
    .A(\memory[4][5] ),
    .B(_01453_),
    .Y(_02869_)
  );
  AND _11035_ (
    .A(_02868_),
    .B(_02869_),
    .Y(_02870_)
  );
  NAND _11036_ (
    .A(\memory[28][5] ),
    .B(_01484_),
    .Y(_02871_)
  );
  NAND _11037_ (
    .A(\memory[7][5] ),
    .B(_01585_),
    .Y(_02872_)
  );
  AND _11038_ (
    .A(_02871_),
    .B(_02872_),
    .Y(_02873_)
  );
  AND _11039_ (
    .A(_02870_),
    .B(_02873_),
    .Y(_02874_)
  );
  NAND _11040_ (
    .A(\memory[2][5] ),
    .B(_01449_),
    .Y(_02875_)
  );
  NAND _11041_ (
    .A(\memory[3][5] ),
    .B(_01570_),
    .Y(_02876_)
  );
  AND _11042_ (
    .A(_02875_),
    .B(_02876_),
    .Y(_02877_)
  );
  NAND _11043_ (
    .A(\memory[16][5] ),
    .B(_01543_),
    .Y(_02878_)
  );
  NAND _11044_ (
    .A(\memory[24][5] ),
    .B(_01469_),
    .Y(_02879_)
  );
  AND _11045_ (
    .A(_02878_),
    .B(_02879_),
    .Y(_02880_)
  );
  AND _11046_ (
    .A(_02877_),
    .B(_02880_),
    .Y(_02881_)
  );
  AND _11047_ (
    .A(_02874_),
    .B(_02881_),
    .Y(_02882_)
  );
  AND _11048_ (
    .A(_02867_),
    .B(_02882_),
    .Y(_02883_)
  );
  NAND _11049_ (
    .A(\memory[25][5] ),
    .B(_01546_),
    .Y(_02884_)
  );
  NAND _11050_ (
    .A(\memory[21][5] ),
    .B(_01534_),
    .Y(_02885_)
  );
  AND _11051_ (
    .A(_02884_),
    .B(_02885_),
    .Y(_02886_)
  );
  NAND _11052_ (
    .A(\memory[11][5] ),
    .B(_01495_),
    .Y(_02887_)
  );
  NAND _11053_ (
    .A(\memory[22][5] ),
    .B(_01553_),
    .Y(_02888_)
  );
  AND _11054_ (
    .A(_02887_),
    .B(_02888_),
    .Y(_02889_)
  );
  AND _11055_ (
    .A(_02886_),
    .B(_02889_),
    .Y(_02890_)
  );
  NAND _11056_ (
    .A(\memory[14][5] ),
    .B(_01458_),
    .Y(_02891_)
  );
  NAND _11057_ (
    .A(\memory[15][5] ),
    .B(_01520_),
    .Y(_02892_)
  );
  AND _11058_ (
    .A(_02891_),
    .B(_02892_),
    .Y(_02893_)
  );
  NAND _11059_ (
    .A(\memory[30][5] ),
    .B(_01462_),
    .Y(_02894_)
  );
  NAND _11060_ (
    .A(\memory[29][5] ),
    .B(_01563_),
    .Y(_02895_)
  );
  AND _11061_ (
    .A(_02894_),
    .B(_02895_),
    .Y(_02896_)
  );
  AND _11062_ (
    .A(_02893_),
    .B(_02896_),
    .Y(_02897_)
  );
  AND _11063_ (
    .A(_02890_),
    .B(_02897_),
    .Y(_02898_)
  );
  NAND _11064_ (
    .A(\memory[17][5] ),
    .B(_01501_),
    .Y(_02899_)
  );
  NAND _11065_ (
    .A(\memory[19][5] ),
    .B(_01479_),
    .Y(_02900_)
  );
  AND _11066_ (
    .A(_02899_),
    .B(_02900_),
    .Y(_02901_)
  );
  NAND _11067_ (
    .A(\memory[0][5] ),
    .B(_01491_),
    .Y(_02902_)
  );
  NAND _11068_ (
    .A(\memory[26][5] ),
    .B(_01550_),
    .Y(_02903_)
  );
  AND _11069_ (
    .A(_02902_),
    .B(_02903_),
    .Y(_02904_)
  );
  AND _11070_ (
    .A(_02901_),
    .B(_02904_),
    .Y(_02905_)
  );
  NAND _11071_ (
    .A(\memory[23][5] ),
    .B(_01474_),
    .Y(_02906_)
  );
  NAND _11072_ (
    .A(\memory[6][5] ),
    .B(_01530_),
    .Y(_02907_)
  );
  AND _11073_ (
    .A(_02906_),
    .B(_02907_),
    .Y(_02908_)
  );
  NAND _11074_ (
    .A(\memory[12][5] ),
    .B(_01578_),
    .Y(_02909_)
  );
  NAND _11075_ (
    .A(\memory[9][5] ),
    .B(_01538_),
    .Y(_02910_)
  );
  AND _11076_ (
    .A(_02909_),
    .B(_02910_),
    .Y(_02911_)
  );
  AND _11077_ (
    .A(_02908_),
    .B(_02911_),
    .Y(_02912_)
  );
  AND _11078_ (
    .A(_02905_),
    .B(_02912_),
    .Y(_02913_)
  );
  AND _11079_ (
    .A(_02898_),
    .B(_02913_),
    .Y(_02914_)
  );
  NAND _11080_ (
    .A(_02883_),
    .B(_02914_),
    .Y(_02915_)
  );
  AND _11081_ (
    .A(MemRead_i),
    .B(_02915_),
    .Y(\data_o[21] )
  );
  NAND _11082_ (
    .A(\memory[5][6] ),
    .B(_01513_),
    .Y(_02916_)
  );
  NAND _11083_ (
    .A(\memory[16][6] ),
    .B(_01543_),
    .Y(_02917_)
  );
  AND _11084_ (
    .A(_02916_),
    .B(_02917_),
    .Y(_02918_)
  );
  NAND _11085_ (
    .A(\memory[23][6] ),
    .B(_01474_),
    .Y(_02919_)
  );
  NAND _11086_ (
    .A(\memory[6][6] ),
    .B(_01530_),
    .Y(_02920_)
  );
  AND _11087_ (
    .A(_02919_),
    .B(_02920_),
    .Y(_02921_)
  );
  AND _11088_ (
    .A(_02918_),
    .B(_02921_),
    .Y(_02922_)
  );
  NAND _11089_ (
    .A(\memory[10][6] ),
    .B(_01527_),
    .Y(_02923_)
  );
  NAND _11090_ (
    .A(\memory[13][6] ),
    .B(_01575_),
    .Y(_02924_)
  );
  AND _11091_ (
    .A(_02923_),
    .B(_02924_),
    .Y(_02925_)
  );
  NAND _11092_ (
    .A(\memory[8][6] ),
    .B(_01517_),
    .Y(_02926_)
  );
  NAND _11093_ (
    .A(\memory[14][6] ),
    .B(_01458_),
    .Y(_02927_)
  );
  AND _11094_ (
    .A(_02926_),
    .B(_02927_),
    .Y(_02928_)
  );
  AND _11095_ (
    .A(_02925_),
    .B(_02928_),
    .Y(_02929_)
  );
  AND _11096_ (
    .A(_02922_),
    .B(_02929_),
    .Y(_02930_)
  );
  NAND _11097_ (
    .A(\memory[3][6] ),
    .B(_01570_),
    .Y(_02931_)
  );
  NAND _11098_ (
    .A(\memory[1][6] ),
    .B(_01504_),
    .Y(_02932_)
  );
  AND _11099_ (
    .A(_02931_),
    .B(_02932_),
    .Y(_02933_)
  );
  NAND _11100_ (
    .A(\memory[19][6] ),
    .B(_01479_),
    .Y(_02934_)
  );
  NAND _11101_ (
    .A(\memory[20][6] ),
    .B(_01582_),
    .Y(_02935_)
  );
  AND _11102_ (
    .A(_02934_),
    .B(_02935_),
    .Y(_02936_)
  );
  AND _11103_ (
    .A(_02933_),
    .B(_02936_),
    .Y(_02937_)
  );
  NAND _11104_ (
    .A(\memory[9][6] ),
    .B(_01538_),
    .Y(_02938_)
  );
  NAND _11105_ (
    .A(\memory[7][6] ),
    .B(_01585_),
    .Y(_02939_)
  );
  AND _11106_ (
    .A(_02938_),
    .B(_02939_),
    .Y(_02940_)
  );
  NAND _11107_ (
    .A(\memory[2][6] ),
    .B(_01449_),
    .Y(_02941_)
  );
  NAND _11108_ (
    .A(\memory[26][6] ),
    .B(_01550_),
    .Y(_02942_)
  );
  AND _11109_ (
    .A(_02941_),
    .B(_02942_),
    .Y(_02943_)
  );
  AND _11110_ (
    .A(_02940_),
    .B(_02943_),
    .Y(_02944_)
  );
  AND _11111_ (
    .A(_02937_),
    .B(_02944_),
    .Y(_02945_)
  );
  AND _11112_ (
    .A(_02930_),
    .B(_02945_),
    .Y(_02946_)
  );
  NAND _11113_ (
    .A(\memory[28][6] ),
    .B(_01484_),
    .Y(_02947_)
  );
  NAND _11114_ (
    .A(\memory[0][6] ),
    .B(_01491_),
    .Y(_02948_)
  );
  AND _11115_ (
    .A(_02947_),
    .B(_02948_),
    .Y(_02949_)
  );
  NAND _11116_ (
    .A(\memory[11][6] ),
    .B(_01495_),
    .Y(_02950_)
  );
  NAND _11117_ (
    .A(\memory[25][6] ),
    .B(_01546_),
    .Y(_02951_)
  );
  AND _11118_ (
    .A(_02950_),
    .B(_02951_),
    .Y(_02952_)
  );
  AND _11119_ (
    .A(_02949_),
    .B(_02952_),
    .Y(_02953_)
  );
  NAND _11120_ (
    .A(\memory[29][6] ),
    .B(_01563_),
    .Y(_02954_)
  );
  NAND _11121_ (
    .A(\memory[31][6] ),
    .B(_01510_),
    .Y(_02955_)
  );
  AND _11122_ (
    .A(_02954_),
    .B(_02955_),
    .Y(_02956_)
  );
  NAND _11123_ (
    .A(\memory[30][6] ),
    .B(_01462_),
    .Y(_02957_)
  );
  NAND _11124_ (
    .A(\memory[27][6] ),
    .B(_01559_),
    .Y(_02958_)
  );
  AND _11125_ (
    .A(_02957_),
    .B(_02958_),
    .Y(_02959_)
  );
  AND _11126_ (
    .A(_02956_),
    .B(_02959_),
    .Y(_02960_)
  );
  AND _11127_ (
    .A(_02953_),
    .B(_02960_),
    .Y(_02961_)
  );
  NAND _11128_ (
    .A(\memory[17][6] ),
    .B(_01501_),
    .Y(_02962_)
  );
  NAND _11129_ (
    .A(\memory[24][6] ),
    .B(_01469_),
    .Y(_02963_)
  );
  AND _11130_ (
    .A(_02962_),
    .B(_02963_),
    .Y(_02964_)
  );
  NAND _11131_ (
    .A(\memory[4][6] ),
    .B(_01453_),
    .Y(_02965_)
  );
  NAND _11132_ (
    .A(\memory[15][6] ),
    .B(_01520_),
    .Y(_02966_)
  );
  AND _11133_ (
    .A(_02965_),
    .B(_02966_),
    .Y(_02967_)
  );
  AND _11134_ (
    .A(_02964_),
    .B(_02967_),
    .Y(_02968_)
  );
  NAND _11135_ (
    .A(\memory[18][6] ),
    .B(_01567_),
    .Y(_02969_)
  );
  NAND _11136_ (
    .A(\memory[22][6] ),
    .B(_01553_),
    .Y(_02970_)
  );
  AND _11137_ (
    .A(_02969_),
    .B(_02970_),
    .Y(_02971_)
  );
  NAND _11138_ (
    .A(\memory[12][6] ),
    .B(_01578_),
    .Y(_02972_)
  );
  NAND _11139_ (
    .A(\memory[21][6] ),
    .B(_01534_),
    .Y(_02973_)
  );
  AND _11140_ (
    .A(_02972_),
    .B(_02973_),
    .Y(_02974_)
  );
  AND _11141_ (
    .A(_02971_),
    .B(_02974_),
    .Y(_02975_)
  );
  AND _11142_ (
    .A(_02968_),
    .B(_02975_),
    .Y(_02976_)
  );
  AND _11143_ (
    .A(_02961_),
    .B(_02976_),
    .Y(_02977_)
  );
  NAND _11144_ (
    .A(_02946_),
    .B(_02977_),
    .Y(_02978_)
  );
  AND _11145_ (
    .A(MemRead_i),
    .B(_02978_),
    .Y(\data_o[22] )
  );
  NAND _11146_ (
    .A(\memory[4][7] ),
    .B(_01453_),
    .Y(_02979_)
  );
  NAND _11147_ (
    .A(\memory[11][7] ),
    .B(_01495_),
    .Y(_02980_)
  );
  AND _11148_ (
    .A(_02979_),
    .B(_02980_),
    .Y(_02981_)
  );
  NAND _11149_ (
    .A(\memory[22][7] ),
    .B(_01553_),
    .Y(_02982_)
  );
  NAND _11150_ (
    .A(\memory[9][7] ),
    .B(_01538_),
    .Y(_02983_)
  );
  AND _11151_ (
    .A(_02982_),
    .B(_02983_),
    .Y(_02984_)
  );
  AND _11152_ (
    .A(_02981_),
    .B(_02984_),
    .Y(_02985_)
  );
  NAND _11153_ (
    .A(\memory[17][7] ),
    .B(_01501_),
    .Y(_02986_)
  );
  NAND _11154_ (
    .A(\memory[3][7] ),
    .B(_01570_),
    .Y(_02987_)
  );
  AND _11155_ (
    .A(_02986_),
    .B(_02987_),
    .Y(_02988_)
  );
  NAND _11156_ (
    .A(\memory[13][7] ),
    .B(_01575_),
    .Y(_02989_)
  );
  NAND _11157_ (
    .A(\memory[15][7] ),
    .B(_01520_),
    .Y(_02990_)
  );
  AND _11158_ (
    .A(_02989_),
    .B(_02990_),
    .Y(_02991_)
  );
  AND _11159_ (
    .A(_02988_),
    .B(_02991_),
    .Y(_02992_)
  );
  AND _11160_ (
    .A(_02985_),
    .B(_02992_),
    .Y(_02993_)
  );
  NAND _11161_ (
    .A(\memory[26][7] ),
    .B(_01550_),
    .Y(_02994_)
  );
  NAND _11162_ (
    .A(\memory[27][7] ),
    .B(_01559_),
    .Y(_02995_)
  );
  AND _11163_ (
    .A(_02994_),
    .B(_02995_),
    .Y(_02996_)
  );
  NAND _11164_ (
    .A(\memory[24][7] ),
    .B(_01469_),
    .Y(_02997_)
  );
  NAND _11165_ (
    .A(\memory[2][7] ),
    .B(_01449_),
    .Y(_02998_)
  );
  AND _11166_ (
    .A(_02997_),
    .B(_02998_),
    .Y(_02999_)
  );
  AND _11167_ (
    .A(_02996_),
    .B(_02999_),
    .Y(_03000_)
  );
  NAND _11168_ (
    .A(\memory[29][7] ),
    .B(_01563_),
    .Y(_03001_)
  );
  NAND _11169_ (
    .A(\memory[31][7] ),
    .B(_01510_),
    .Y(_03002_)
  );
  AND _11170_ (
    .A(_03001_),
    .B(_03002_),
    .Y(_03003_)
  );
  NAND _11171_ (
    .A(\memory[19][7] ),
    .B(_01479_),
    .Y(_03004_)
  );
  NAND _11172_ (
    .A(\memory[21][7] ),
    .B(_01534_),
    .Y(_03005_)
  );
  AND _11173_ (
    .A(_03004_),
    .B(_03005_),
    .Y(_03006_)
  );
  AND _11174_ (
    .A(_03003_),
    .B(_03006_),
    .Y(_03007_)
  );
  AND _11175_ (
    .A(_03000_),
    .B(_03007_),
    .Y(_03008_)
  );
  AND _11176_ (
    .A(_02993_),
    .B(_03008_),
    .Y(_03009_)
  );
  NAND _11177_ (
    .A(\memory[6][7] ),
    .B(_01530_),
    .Y(_03010_)
  );
  NAND _11178_ (
    .A(\memory[8][7] ),
    .B(_01517_),
    .Y(_03011_)
  );
  AND _11179_ (
    .A(_03010_),
    .B(_03011_),
    .Y(_03012_)
  );
  NAND _11180_ (
    .A(\memory[5][7] ),
    .B(_01513_),
    .Y(_03013_)
  );
  NAND _11181_ (
    .A(\memory[28][7] ),
    .B(_01484_),
    .Y(_03014_)
  );
  AND _11182_ (
    .A(_03013_),
    .B(_03014_),
    .Y(_03015_)
  );
  AND _11183_ (
    .A(_03012_),
    .B(_03015_),
    .Y(_03016_)
  );
  NAND _11184_ (
    .A(\memory[10][7] ),
    .B(_01527_),
    .Y(_03017_)
  );
  NAND _11185_ (
    .A(\memory[14][7] ),
    .B(_01458_),
    .Y(_03018_)
  );
  AND _11186_ (
    .A(_03017_),
    .B(_03018_),
    .Y(_03019_)
  );
  NAND _11187_ (
    .A(\memory[25][7] ),
    .B(_01546_),
    .Y(_03020_)
  );
  NAND _11188_ (
    .A(\memory[20][7] ),
    .B(_01582_),
    .Y(_03021_)
  );
  AND _11189_ (
    .A(_03020_),
    .B(_03021_),
    .Y(_03022_)
  );
  AND _11190_ (
    .A(_03019_),
    .B(_03022_),
    .Y(_03023_)
  );
  AND _11191_ (
    .A(_03016_),
    .B(_03023_),
    .Y(_03024_)
  );
  NAND _11192_ (
    .A(\memory[12][7] ),
    .B(_01578_),
    .Y(_03025_)
  );
  NAND _11193_ (
    .A(\memory[16][7] ),
    .B(_01543_),
    .Y(_03026_)
  );
  AND _11194_ (
    .A(_03025_),
    .B(_03026_),
    .Y(_03027_)
  );
  NAND _11195_ (
    .A(\memory[7][7] ),
    .B(_01585_),
    .Y(_03028_)
  );
  NAND _11196_ (
    .A(\memory[1][7] ),
    .B(_01504_),
    .Y(_03029_)
  );
  AND _11197_ (
    .A(_03028_),
    .B(_03029_),
    .Y(_03030_)
  );
  AND _11198_ (
    .A(_03027_),
    .B(_03030_),
    .Y(_03031_)
  );
  NAND _11199_ (
    .A(\memory[23][7] ),
    .B(_01474_),
    .Y(_03032_)
  );
  NAND _11200_ (
    .A(\memory[30][7] ),
    .B(_01462_),
    .Y(_03033_)
  );
  AND _11201_ (
    .A(_03032_),
    .B(_03033_),
    .Y(_03034_)
  );
  NAND _11202_ (
    .A(\memory[18][7] ),
    .B(_01567_),
    .Y(_03035_)
  );
  NAND _11203_ (
    .A(\memory[0][7] ),
    .B(_01491_),
    .Y(_03036_)
  );
  AND _11204_ (
    .A(_03035_),
    .B(_03036_),
    .Y(_03037_)
  );
  AND _11205_ (
    .A(_03034_),
    .B(_03037_),
    .Y(_03038_)
  );
  AND _11206_ (
    .A(_03031_),
    .B(_03038_),
    .Y(_03039_)
  );
  AND _11207_ (
    .A(_03024_),
    .B(_03039_),
    .Y(_03040_)
  );
  NAND _11208_ (
    .A(_03009_),
    .B(_03040_),
    .Y(_03041_)
  );
  AND _11209_ (
    .A(MemRead_i),
    .B(_03041_),
    .Y(\data_o[23] )
  );
  NAND _11210_ (
    .A(\memory[20][0] ),
    .B(_01479_),
    .Y(_03042_)
  );
  NAND _11211_ (
    .A(\memory[9][0] ),
    .B(_01517_),
    .Y(_03043_)
  );
  AND _11212_ (
    .A(_03042_),
    .B(_03043_),
    .Y(_03044_)
  );
  NAND _11213_ (
    .A(\memory[6][0] ),
    .B(_01513_),
    .Y(_03045_)
  );
  NAND _11214_ (
    .A(\memory[4][0] ),
    .B(_01570_),
    .Y(_03046_)
  );
  AND _11215_ (
    .A(_03045_),
    .B(_03046_),
    .Y(_03047_)
  );
  AND _11216_ (
    .A(_03044_),
    .B(_03047_),
    .Y(_03048_)
  );
  NAND _11217_ (
    .A(\memory[16][0] ),
    .B(_01520_),
    .Y(_03049_)
  );
  NAND _11218_ (
    .A(\memory[3][0] ),
    .B(_01449_),
    .Y(_03050_)
  );
  AND _11219_ (
    .A(_03049_),
    .B(_03050_),
    .Y(_03051_)
  );
  NAND _11220_ (
    .A(\memory[25][0] ),
    .B(_01469_),
    .Y(_03052_)
  );
  NAND _11221_ (
    .A(\memory[15][0] ),
    .B(_01458_),
    .Y(_03053_)
  );
  AND _11222_ (
    .A(_03052_),
    .B(_03053_),
    .Y(_03054_)
  );
  AND _11223_ (
    .A(_03051_),
    .B(_03054_),
    .Y(_03055_)
  );
  AND _11224_ (
    .A(_03048_),
    .B(_03055_),
    .Y(_03056_)
  );
  NAND _11225_ (
    .A(\memory[28][0] ),
    .B(_01559_),
    .Y(_03057_)
  );
  NAND _11226_ (
    .A(\memory[22][0] ),
    .B(_01534_),
    .Y(_03058_)
  );
  AND _11227_ (
    .A(_03057_),
    .B(_03058_),
    .Y(_03059_)
  );
  NAND _11228_ (
    .A(\memory[8][0] ),
    .B(_01585_),
    .Y(_03060_)
  );
  NAND _11229_ (
    .A(\memory[0][0] ),
    .B(_01510_),
    .Y(_03061_)
  );
  AND _11230_ (
    .A(_03060_),
    .B(_03061_),
    .Y(_03062_)
  );
  AND _11231_ (
    .A(_03059_),
    .B(_03062_),
    .Y(_03063_)
  );
  NAND _11232_ (
    .A(\memory[7][0] ),
    .B(_01530_),
    .Y(_03064_)
  );
  NAND _11233_ (
    .A(\memory[24][0] ),
    .B(_01474_),
    .Y(_03065_)
  );
  AND _11234_ (
    .A(_03064_),
    .B(_03065_),
    .Y(_03066_)
  );
  NAND _11235_ (
    .A(\memory[18][0] ),
    .B(_01501_),
    .Y(_03067_)
  );
  NAND _11236_ (
    .A(\memory[5][0] ),
    .B(_01453_),
    .Y(_03068_)
  );
  AND _11237_ (
    .A(_03067_),
    .B(_03068_),
    .Y(_03069_)
  );
  AND _11238_ (
    .A(_03066_),
    .B(_03069_),
    .Y(_03070_)
  );
  AND _11239_ (
    .A(_03063_),
    .B(_03070_),
    .Y(_03071_)
  );
  AND _11240_ (
    .A(_03056_),
    .B(_03071_),
    .Y(_03072_)
  );
  NAND _11241_ (
    .A(\memory[2][0] ),
    .B(_01504_),
    .Y(_03073_)
  );
  NAND _11242_ (
    .A(\memory[1][0] ),
    .B(_01491_),
    .Y(_03074_)
  );
  AND _11243_ (
    .A(_03073_),
    .B(_03074_),
    .Y(_03075_)
  );
  NAND _11244_ (
    .A(\memory[21][0] ),
    .B(_01582_),
    .Y(_03076_)
  );
  NAND _11245_ (
    .A(\memory[12][0] ),
    .B(_01495_),
    .Y(_03077_)
  );
  AND _11246_ (
    .A(_03076_),
    .B(_03077_),
    .Y(_03078_)
  );
  AND _11247_ (
    .A(_03075_),
    .B(_03078_),
    .Y(_03079_)
  );
  NAND _11248_ (
    .A(\memory[14][0] ),
    .B(_01575_),
    .Y(_03080_)
  );
  NAND _11249_ (
    .A(\memory[30][0] ),
    .B(_01563_),
    .Y(_03081_)
  );
  AND _11250_ (
    .A(_03080_),
    .B(_03081_),
    .Y(_03082_)
  );
  NAND _11251_ (
    .A(\memory[27][0] ),
    .B(_01550_),
    .Y(_03083_)
  );
  NAND _11252_ (
    .A(\memory[29][0] ),
    .B(_01484_),
    .Y(_03084_)
  );
  AND _11253_ (
    .A(_03083_),
    .B(_03084_),
    .Y(_03085_)
  );
  AND _11254_ (
    .A(_03082_),
    .B(_03085_),
    .Y(_03086_)
  );
  AND _11255_ (
    .A(_03079_),
    .B(_03086_),
    .Y(_03087_)
  );
  NAND _11256_ (
    .A(\memory[11][0] ),
    .B(_01527_),
    .Y(_03088_)
  );
  NAND _11257_ (
    .A(\memory[10][0] ),
    .B(_01538_),
    .Y(_03089_)
  );
  AND _11258_ (
    .A(_03088_),
    .B(_03089_),
    .Y(_03090_)
  );
  NAND _11259_ (
    .A(\memory[19][0] ),
    .B(_01567_),
    .Y(_03091_)
  );
  NAND _11260_ (
    .A(\memory[23][0] ),
    .B(_01553_),
    .Y(_03092_)
  );
  AND _11261_ (
    .A(_03091_),
    .B(_03092_),
    .Y(_03093_)
  );
  AND _11262_ (
    .A(_03090_),
    .B(_03093_),
    .Y(_03094_)
  );
  NAND _11263_ (
    .A(\memory[17][0] ),
    .B(_01543_),
    .Y(_03095_)
  );
  NAND _11264_ (
    .A(\memory[26][0] ),
    .B(_01546_),
    .Y(_03096_)
  );
  AND _11265_ (
    .A(_03095_),
    .B(_03096_),
    .Y(_03097_)
  );
  NAND _11266_ (
    .A(\memory[31][0] ),
    .B(_01462_),
    .Y(_03098_)
  );
  NAND _11267_ (
    .A(\memory[13][0] ),
    .B(_01578_),
    .Y(_03099_)
  );
  AND _11268_ (
    .A(_03098_),
    .B(_03099_),
    .Y(_03100_)
  );
  AND _11269_ (
    .A(_03097_),
    .B(_03100_),
    .Y(_03101_)
  );
  AND _11270_ (
    .A(_03094_),
    .B(_03101_),
    .Y(_03102_)
  );
  AND _11271_ (
    .A(_03087_),
    .B(_03102_),
    .Y(_03103_)
  );
  NAND _11272_ (
    .A(_03072_),
    .B(_03103_),
    .Y(_03104_)
  );
  AND _11273_ (
    .A(MemRead_i),
    .B(_03104_),
    .Y(\data_o[24] )
  );
  NAND _11274_ (
    .A(\memory[13][1] ),
    .B(_01578_),
    .Y(_03105_)
  );
  NAND _11275_ (
    .A(\memory[11][1] ),
    .B(_01527_),
    .Y(_03106_)
  );
  AND _11276_ (
    .A(_03105_),
    .B(_03106_),
    .Y(_03107_)
  );
  NAND _11277_ (
    .A(\memory[24][1] ),
    .B(_01474_),
    .Y(_03108_)
  );
  NAND _11278_ (
    .A(\memory[6][1] ),
    .B(_01513_),
    .Y(_03109_)
  );
  AND _11279_ (
    .A(_03108_),
    .B(_03109_),
    .Y(_03110_)
  );
  AND _11280_ (
    .A(_03107_),
    .B(_03110_),
    .Y(_03111_)
  );
  NAND _11281_ (
    .A(\memory[28][1] ),
    .B(_01559_),
    .Y(_03112_)
  );
  NAND _11282_ (
    .A(\memory[8][1] ),
    .B(_01585_),
    .Y(_03113_)
  );
  AND _11283_ (
    .A(_03112_),
    .B(_03113_),
    .Y(_03114_)
  );
  NAND _11284_ (
    .A(\memory[10][1] ),
    .B(_01538_),
    .Y(_03115_)
  );
  NAND _11285_ (
    .A(\memory[18][1] ),
    .B(_01501_),
    .Y(_03116_)
  );
  AND _11286_ (
    .A(_03115_),
    .B(_03116_),
    .Y(_03117_)
  );
  AND _11287_ (
    .A(_03114_),
    .B(_03117_),
    .Y(_03118_)
  );
  AND _11288_ (
    .A(_03111_),
    .B(_03118_),
    .Y(_03119_)
  );
  NAND _11289_ (
    .A(\memory[30][1] ),
    .B(_01563_),
    .Y(_03120_)
  );
  NAND _11290_ (
    .A(\memory[0][1] ),
    .B(_01510_),
    .Y(_03121_)
  );
  AND _11291_ (
    .A(_03120_),
    .B(_03121_),
    .Y(_03122_)
  );
  NAND _11292_ (
    .A(\memory[31][1] ),
    .B(_01462_),
    .Y(_03123_)
  );
  NAND _11293_ (
    .A(\memory[25][1] ),
    .B(_01469_),
    .Y(_03124_)
  );
  AND _11294_ (
    .A(_03123_),
    .B(_03124_),
    .Y(_03125_)
  );
  AND _11295_ (
    .A(_03122_),
    .B(_03125_),
    .Y(_03126_)
  );
  NAND _11296_ (
    .A(\memory[4][1] ),
    .B(_01570_),
    .Y(_03127_)
  );
  NAND _11297_ (
    .A(\memory[7][1] ),
    .B(_01530_),
    .Y(_03128_)
  );
  AND _11298_ (
    .A(_03127_),
    .B(_03128_),
    .Y(_03129_)
  );
  NAND _11299_ (
    .A(\memory[20][1] ),
    .B(_01479_),
    .Y(_03130_)
  );
  NAND _11300_ (
    .A(\memory[26][1] ),
    .B(_01546_),
    .Y(_03131_)
  );
  AND _11301_ (
    .A(_03130_),
    .B(_03131_),
    .Y(_03132_)
  );
  AND _11302_ (
    .A(_03129_),
    .B(_03132_),
    .Y(_03133_)
  );
  AND _11303_ (
    .A(_03126_),
    .B(_03133_),
    .Y(_03134_)
  );
  AND _11304_ (
    .A(_03119_),
    .B(_03134_),
    .Y(_03135_)
  );
  NAND _11305_ (
    .A(\memory[16][1] ),
    .B(_01520_),
    .Y(_03136_)
  );
  NAND _11306_ (
    .A(\memory[19][1] ),
    .B(_01567_),
    .Y(_03137_)
  );
  AND _11307_ (
    .A(_03136_),
    .B(_03137_),
    .Y(_03138_)
  );
  NAND _11308_ (
    .A(\memory[9][1] ),
    .B(_01517_),
    .Y(_03139_)
  );
  NAND _11309_ (
    .A(\memory[5][1] ),
    .B(_01453_),
    .Y(_03140_)
  );
  AND _11310_ (
    .A(_03139_),
    .B(_03140_),
    .Y(_03141_)
  );
  AND _11311_ (
    .A(_03138_),
    .B(_03141_),
    .Y(_03142_)
  );
  NAND _11312_ (
    .A(\memory[22][1] ),
    .B(_01534_),
    .Y(_03143_)
  );
  NAND _11313_ (
    .A(\memory[12][1] ),
    .B(_01495_),
    .Y(_03144_)
  );
  AND _11314_ (
    .A(_03143_),
    .B(_03144_),
    .Y(_03145_)
  );
  NAND _11315_ (
    .A(\memory[17][1] ),
    .B(_01543_),
    .Y(_03146_)
  );
  NAND _11316_ (
    .A(\memory[1][1] ),
    .B(_01491_),
    .Y(_03147_)
  );
  AND _11317_ (
    .A(_03146_),
    .B(_03147_),
    .Y(_03148_)
  );
  AND _11318_ (
    .A(_03145_),
    .B(_03148_),
    .Y(_03149_)
  );
  AND _11319_ (
    .A(_03142_),
    .B(_03149_),
    .Y(_03150_)
  );
  NAND _11320_ (
    .A(\memory[29][1] ),
    .B(_01484_),
    .Y(_03151_)
  );
  NAND _11321_ (
    .A(\memory[14][1] ),
    .B(_01575_),
    .Y(_03152_)
  );
  AND _11322_ (
    .A(_03151_),
    .B(_03152_),
    .Y(_03153_)
  );
  NAND _11323_ (
    .A(\memory[27][1] ),
    .B(_01550_),
    .Y(_03154_)
  );
  NAND _11324_ (
    .A(\memory[23][1] ),
    .B(_01553_),
    .Y(_03155_)
  );
  AND _11325_ (
    .A(_03154_),
    .B(_03155_),
    .Y(_03156_)
  );
  AND _11326_ (
    .A(_03153_),
    .B(_03156_),
    .Y(_03157_)
  );
  NAND _11327_ (
    .A(\memory[21][1] ),
    .B(_01582_),
    .Y(_03158_)
  );
  NAND _11328_ (
    .A(\memory[15][1] ),
    .B(_01458_),
    .Y(_03159_)
  );
  AND _11329_ (
    .A(_03158_),
    .B(_03159_),
    .Y(_03160_)
  );
  NAND _11330_ (
    .A(\memory[3][1] ),
    .B(_01449_),
    .Y(_03161_)
  );
  NAND _11331_ (
    .A(\memory[2][1] ),
    .B(_01504_),
    .Y(_03162_)
  );
  AND _11332_ (
    .A(_03161_),
    .B(_03162_),
    .Y(_03163_)
  );
  AND _11333_ (
    .A(_03160_),
    .B(_03163_),
    .Y(_03164_)
  );
  AND _11334_ (
    .A(_03157_),
    .B(_03164_),
    .Y(_03165_)
  );
  AND _11335_ (
    .A(_03150_),
    .B(_03165_),
    .Y(_03166_)
  );
  NAND _11336_ (
    .A(_03135_),
    .B(_03166_),
    .Y(_03167_)
  );
  AND _11337_ (
    .A(MemRead_i),
    .B(_03167_),
    .Y(\data_o[25] )
  );
  NAND _11338_ (
    .A(\memory[24][2] ),
    .B(_01474_),
    .Y(_03168_)
  );
  NAND _11339_ (
    .A(\memory[30][2] ),
    .B(_01563_),
    .Y(_03169_)
  );
  AND _11340_ (
    .A(_03168_),
    .B(_03169_),
    .Y(_03170_)
  );
  NAND _11341_ (
    .A(\memory[8][2] ),
    .B(_01585_),
    .Y(_03171_)
  );
  NAND _11342_ (
    .A(\memory[15][2] ),
    .B(_01458_),
    .Y(_03172_)
  );
  AND _11343_ (
    .A(_03171_),
    .B(_03172_),
    .Y(_03173_)
  );
  AND _11344_ (
    .A(_03170_),
    .B(_03173_),
    .Y(_03174_)
  );
  NAND _11345_ (
    .A(\memory[28][2] ),
    .B(_01559_),
    .Y(_03175_)
  );
  NAND _11346_ (
    .A(\memory[5][2] ),
    .B(_01453_),
    .Y(_03176_)
  );
  AND _11347_ (
    .A(_03175_),
    .B(_03176_),
    .Y(_03177_)
  );
  NAND _11348_ (
    .A(\memory[22][2] ),
    .B(_01534_),
    .Y(_03178_)
  );
  NAND _11349_ (
    .A(\memory[23][2] ),
    .B(_01553_),
    .Y(_03179_)
  );
  AND _11350_ (
    .A(_03178_),
    .B(_03179_),
    .Y(_03180_)
  );
  AND _11351_ (
    .A(_03177_),
    .B(_03180_),
    .Y(_03181_)
  );
  AND _11352_ (
    .A(_03174_),
    .B(_03181_),
    .Y(_03182_)
  );
  NAND _11353_ (
    .A(\memory[17][2] ),
    .B(_01543_),
    .Y(_03183_)
  );
  NAND _11354_ (
    .A(\memory[20][2] ),
    .B(_01479_),
    .Y(_03184_)
  );
  AND _11355_ (
    .A(_03183_),
    .B(_03184_),
    .Y(_03185_)
  );
  NAND _11356_ (
    .A(\memory[3][2] ),
    .B(_01449_),
    .Y(_03186_)
  );
  NAND _11357_ (
    .A(\memory[1][2] ),
    .B(_01491_),
    .Y(_03187_)
  );
  AND _11358_ (
    .A(_03186_),
    .B(_03187_),
    .Y(_03188_)
  );
  AND _11359_ (
    .A(_03185_),
    .B(_03188_),
    .Y(_03189_)
  );
  NAND _11360_ (
    .A(\memory[18][2] ),
    .B(_01501_),
    .Y(_03190_)
  );
  NAND _11361_ (
    .A(\memory[19][2] ),
    .B(_01567_),
    .Y(_03191_)
  );
  AND _11362_ (
    .A(_03190_),
    .B(_03191_),
    .Y(_03192_)
  );
  NAND _11363_ (
    .A(\memory[7][2] ),
    .B(_01530_),
    .Y(_03193_)
  );
  NAND _11364_ (
    .A(\memory[14][2] ),
    .B(_01575_),
    .Y(_03194_)
  );
  AND _11365_ (
    .A(_03193_),
    .B(_03194_),
    .Y(_03195_)
  );
  AND _11366_ (
    .A(_03192_),
    .B(_03195_),
    .Y(_03196_)
  );
  AND _11367_ (
    .A(_03189_),
    .B(_03196_),
    .Y(_03197_)
  );
  AND _11368_ (
    .A(_03182_),
    .B(_03197_),
    .Y(_03198_)
  );
  NAND _11369_ (
    .A(\memory[27][2] ),
    .B(_01550_),
    .Y(_03199_)
  );
  NAND _11370_ (
    .A(\memory[31][2] ),
    .B(_01462_),
    .Y(_03200_)
  );
  AND _11371_ (
    .A(_03199_),
    .B(_03200_),
    .Y(_03201_)
  );
  NAND _11372_ (
    .A(\memory[26][2] ),
    .B(_01546_),
    .Y(_03202_)
  );
  NAND _11373_ (
    .A(\memory[12][2] ),
    .B(_01495_),
    .Y(_03203_)
  );
  AND _11374_ (
    .A(_03202_),
    .B(_03203_),
    .Y(_03204_)
  );
  AND _11375_ (
    .A(_03201_),
    .B(_03204_),
    .Y(_03205_)
  );
  NAND _11376_ (
    .A(\memory[25][2] ),
    .B(_01469_),
    .Y(_03206_)
  );
  NAND _11377_ (
    .A(\memory[4][2] ),
    .B(_01570_),
    .Y(_03207_)
  );
  AND _11378_ (
    .A(_03206_),
    .B(_03207_),
    .Y(_03208_)
  );
  NAND _11379_ (
    .A(\memory[16][2] ),
    .B(_01520_),
    .Y(_03209_)
  );
  NAND _11380_ (
    .A(\memory[13][2] ),
    .B(_01578_),
    .Y(_03210_)
  );
  AND _11381_ (
    .A(_03209_),
    .B(_03210_),
    .Y(_03211_)
  );
  AND _11382_ (
    .A(_03208_),
    .B(_03211_),
    .Y(_03212_)
  );
  AND _11383_ (
    .A(_03205_),
    .B(_03212_),
    .Y(_03213_)
  );
  NAND _11384_ (
    .A(\memory[10][2] ),
    .B(_01538_),
    .Y(_03214_)
  );
  NAND _11385_ (
    .A(\memory[11][2] ),
    .B(_01527_),
    .Y(_03215_)
  );
  AND _11386_ (
    .A(_03214_),
    .B(_03215_),
    .Y(_03216_)
  );
  NAND _11387_ (
    .A(\memory[2][2] ),
    .B(_01504_),
    .Y(_03217_)
  );
  NAND _11388_ (
    .A(\memory[0][2] ),
    .B(_01510_),
    .Y(_03218_)
  );
  AND _11389_ (
    .A(_03217_),
    .B(_03218_),
    .Y(_03219_)
  );
  AND _11390_ (
    .A(_03216_),
    .B(_03219_),
    .Y(_03220_)
  );
  NAND _11391_ (
    .A(\memory[6][2] ),
    .B(_01513_),
    .Y(_03221_)
  );
  NAND _11392_ (
    .A(\memory[9][2] ),
    .B(_01517_),
    .Y(_03222_)
  );
  AND _11393_ (
    .A(_03221_),
    .B(_03222_),
    .Y(_03223_)
  );
  NAND _11394_ (
    .A(\memory[29][2] ),
    .B(_01484_),
    .Y(_03224_)
  );
  NAND _11395_ (
    .A(\memory[21][2] ),
    .B(_01582_),
    .Y(_03225_)
  );
  AND _11396_ (
    .A(_03224_),
    .B(_03225_),
    .Y(_03226_)
  );
  AND _11397_ (
    .A(_03223_),
    .B(_03226_),
    .Y(_03227_)
  );
  AND _11398_ (
    .A(_03220_),
    .B(_03227_),
    .Y(_03228_)
  );
  AND _11399_ (
    .A(_03213_),
    .B(_03228_),
    .Y(_03229_)
  );
  NAND _11400_ (
    .A(_03198_),
    .B(_03229_),
    .Y(_03230_)
  );
  AND _11401_ (
    .A(MemRead_i),
    .B(_03230_),
    .Y(\data_o[26] )
  );
  NAND _11402_ (
    .A(\memory[13][3] ),
    .B(_01578_),
    .Y(_03231_)
  );
  NAND _11403_ (
    .A(\memory[7][3] ),
    .B(_01530_),
    .Y(_03232_)
  );
  AND _11404_ (
    .A(_03231_),
    .B(_03232_),
    .Y(_03233_)
  );
  NAND _11405_ (
    .A(\memory[14][3] ),
    .B(_01575_),
    .Y(_03234_)
  );
  NAND _11406_ (
    .A(\memory[26][3] ),
    .B(_01546_),
    .Y(_03235_)
  );
  AND _11407_ (
    .A(_03234_),
    .B(_03235_),
    .Y(_03236_)
  );
  AND _11408_ (
    .A(_03233_),
    .B(_03236_),
    .Y(_03237_)
  );
  NAND _11409_ (
    .A(\memory[16][3] ),
    .B(_01520_),
    .Y(_03238_)
  );
  NAND _11410_ (
    .A(\memory[6][3] ),
    .B(_01513_),
    .Y(_03239_)
  );
  AND _11411_ (
    .A(_03238_),
    .B(_03239_),
    .Y(_03240_)
  );
  NAND _11412_ (
    .A(\memory[17][3] ),
    .B(_01543_),
    .Y(_03241_)
  );
  NAND _11413_ (
    .A(\memory[5][3] ),
    .B(_01453_),
    .Y(_03242_)
  );
  AND _11414_ (
    .A(_03241_),
    .B(_03242_),
    .Y(_03243_)
  );
  AND _11415_ (
    .A(_03240_),
    .B(_03243_),
    .Y(_03244_)
  );
  AND _11416_ (
    .A(_03237_),
    .B(_03244_),
    .Y(_03245_)
  );
  NAND _11417_ (
    .A(\memory[0][3] ),
    .B(_01510_),
    .Y(_03246_)
  );
  NAND _11418_ (
    .A(\memory[30][3] ),
    .B(_01563_),
    .Y(_03247_)
  );
  AND _11419_ (
    .A(_03246_),
    .B(_03247_),
    .Y(_03248_)
  );
  NAND _11420_ (
    .A(\memory[11][3] ),
    .B(_01527_),
    .Y(_03249_)
  );
  NAND _11421_ (
    .A(\memory[31][3] ),
    .B(_01462_),
    .Y(_03250_)
  );
  AND _11422_ (
    .A(_03249_),
    .B(_03250_),
    .Y(_03251_)
  );
  AND _11423_ (
    .A(_03248_),
    .B(_03251_),
    .Y(_03252_)
  );
  NAND _11424_ (
    .A(\memory[10][3] ),
    .B(_01538_),
    .Y(_03253_)
  );
  NAND _11425_ (
    .A(\memory[27][3] ),
    .B(_01550_),
    .Y(_03254_)
  );
  AND _11426_ (
    .A(_03253_),
    .B(_03254_),
    .Y(_03255_)
  );
  NAND _11427_ (
    .A(\memory[24][3] ),
    .B(_01474_),
    .Y(_03256_)
  );
  NAND _11428_ (
    .A(\memory[20][3] ),
    .B(_01479_),
    .Y(_03257_)
  );
  AND _11429_ (
    .A(_03256_),
    .B(_03257_),
    .Y(_03258_)
  );
  AND _11430_ (
    .A(_03255_),
    .B(_03258_),
    .Y(_03259_)
  );
  AND _11431_ (
    .A(_03252_),
    .B(_03259_),
    .Y(_03260_)
  );
  AND _11432_ (
    .A(_03245_),
    .B(_03260_),
    .Y(_03261_)
  );
  NAND _11433_ (
    .A(\memory[25][3] ),
    .B(_01469_),
    .Y(_03262_)
  );
  NAND _11434_ (
    .A(\memory[23][3] ),
    .B(_01553_),
    .Y(_03263_)
  );
  AND _11435_ (
    .A(_03262_),
    .B(_03263_),
    .Y(_03264_)
  );
  NAND _11436_ (
    .A(\memory[29][3] ),
    .B(_01484_),
    .Y(_03265_)
  );
  NAND _11437_ (
    .A(\memory[18][3] ),
    .B(_01501_),
    .Y(_03266_)
  );
  AND _11438_ (
    .A(_03265_),
    .B(_03266_),
    .Y(_03267_)
  );
  AND _11439_ (
    .A(_03264_),
    .B(_03267_),
    .Y(_03268_)
  );
  NAND _11440_ (
    .A(\memory[12][3] ),
    .B(_01495_),
    .Y(_03269_)
  );
  NAND _11441_ (
    .A(\memory[15][3] ),
    .B(_01458_),
    .Y(_03270_)
  );
  AND _11442_ (
    .A(_03269_),
    .B(_03270_),
    .Y(_03271_)
  );
  NAND _11443_ (
    .A(\memory[21][3] ),
    .B(_01582_),
    .Y(_03272_)
  );
  NAND _11444_ (
    .A(\memory[22][3] ),
    .B(_01534_),
    .Y(_03273_)
  );
  AND _11445_ (
    .A(_03272_),
    .B(_03273_),
    .Y(_03274_)
  );
  AND _11446_ (
    .A(_03271_),
    .B(_03274_),
    .Y(_03275_)
  );
  AND _11447_ (
    .A(_03268_),
    .B(_03275_),
    .Y(_03276_)
  );
  NAND _11448_ (
    .A(\memory[3][3] ),
    .B(_01449_),
    .Y(_03277_)
  );
  NAND _11449_ (
    .A(\memory[1][3] ),
    .B(_01491_),
    .Y(_03278_)
  );
  AND _11450_ (
    .A(_03277_),
    .B(_03278_),
    .Y(_03279_)
  );
  NAND _11451_ (
    .A(\memory[2][3] ),
    .B(_01504_),
    .Y(_03280_)
  );
  NAND _11452_ (
    .A(\memory[9][3] ),
    .B(_01517_),
    .Y(_03281_)
  );
  AND _11453_ (
    .A(_03280_),
    .B(_03281_),
    .Y(_03282_)
  );
  AND _11454_ (
    .A(_03279_),
    .B(_03282_),
    .Y(_03283_)
  );
  NAND _11455_ (
    .A(\memory[4][3] ),
    .B(_01570_),
    .Y(_03284_)
  );
  NAND _11456_ (
    .A(\memory[19][3] ),
    .B(_01567_),
    .Y(_03285_)
  );
  AND _11457_ (
    .A(_03284_),
    .B(_03285_),
    .Y(_03286_)
  );
  NAND _11458_ (
    .A(\memory[28][3] ),
    .B(_01559_),
    .Y(_03287_)
  );
  NAND _11459_ (
    .A(\memory[8][3] ),
    .B(_01585_),
    .Y(_03288_)
  );
  AND _11460_ (
    .A(_03287_),
    .B(_03288_),
    .Y(_03289_)
  );
  AND _11461_ (
    .A(_03286_),
    .B(_03289_),
    .Y(_03290_)
  );
  AND _11462_ (
    .A(_03283_),
    .B(_03290_),
    .Y(_03291_)
  );
  AND _11463_ (
    .A(_03276_),
    .B(_03291_),
    .Y(_03292_)
  );
  NAND _11464_ (
    .A(_03261_),
    .B(_03292_),
    .Y(_03293_)
  );
  AND _11465_ (
    .A(MemRead_i),
    .B(_03293_),
    .Y(\data_o[27] )
  );
  NAND _11466_ (
    .A(\memory[17][4] ),
    .B(_01543_),
    .Y(_03294_)
  );
  NAND _11467_ (
    .A(\memory[11][4] ),
    .B(_01527_),
    .Y(_03295_)
  );
  AND _11468_ (
    .A(_03294_),
    .B(_03295_),
    .Y(_03296_)
  );
  NAND _11469_ (
    .A(\memory[21][4] ),
    .B(_01582_),
    .Y(_03297_)
  );
  NAND _11470_ (
    .A(\memory[29][4] ),
    .B(_01484_),
    .Y(_03298_)
  );
  AND _11471_ (
    .A(_03297_),
    .B(_03298_),
    .Y(_03299_)
  );
  AND _11472_ (
    .A(_03296_),
    .B(_03299_),
    .Y(_03300_)
  );
  NAND _11473_ (
    .A(\memory[7][4] ),
    .B(_01530_),
    .Y(_03301_)
  );
  NAND _11474_ (
    .A(\memory[1][4] ),
    .B(_01491_),
    .Y(_03302_)
  );
  AND _11475_ (
    .A(_03301_),
    .B(_03302_),
    .Y(_03303_)
  );
  NAND _11476_ (
    .A(\memory[30][4] ),
    .B(_01563_),
    .Y(_03304_)
  );
  NAND _11477_ (
    .A(\memory[28][4] ),
    .B(_01559_),
    .Y(_03305_)
  );
  AND _11478_ (
    .A(_03304_),
    .B(_03305_),
    .Y(_03306_)
  );
  AND _11479_ (
    .A(_03303_),
    .B(_03306_),
    .Y(_03307_)
  );
  AND _11480_ (
    .A(_03300_),
    .B(_03307_),
    .Y(_03308_)
  );
  NAND _11481_ (
    .A(\memory[18][4] ),
    .B(_01501_),
    .Y(_03309_)
  );
  NAND _11482_ (
    .A(\memory[10][4] ),
    .B(_01538_),
    .Y(_03310_)
  );
  AND _11483_ (
    .A(_03309_),
    .B(_03310_),
    .Y(_03311_)
  );
  NAND _11484_ (
    .A(\memory[19][4] ),
    .B(_01567_),
    .Y(_03312_)
  );
  NAND _11485_ (
    .A(\memory[12][4] ),
    .B(_01495_),
    .Y(_03313_)
  );
  AND _11486_ (
    .A(_03312_),
    .B(_03313_),
    .Y(_03314_)
  );
  AND _11487_ (
    .A(_03311_),
    .B(_03314_),
    .Y(_03315_)
  );
  NAND _11488_ (
    .A(\memory[23][4] ),
    .B(_01553_),
    .Y(_03316_)
  );
  NAND _11489_ (
    .A(\memory[14][4] ),
    .B(_01575_),
    .Y(_03317_)
  );
  AND _11490_ (
    .A(_03316_),
    .B(_03317_),
    .Y(_03318_)
  );
  NAND _11491_ (
    .A(\memory[22][4] ),
    .B(_01534_),
    .Y(_03319_)
  );
  NAND _11492_ (
    .A(\memory[0][4] ),
    .B(_01510_),
    .Y(_03320_)
  );
  AND _11493_ (
    .A(_03319_),
    .B(_03320_),
    .Y(_03321_)
  );
  AND _11494_ (
    .A(_03318_),
    .B(_03321_),
    .Y(_03322_)
  );
  AND _11495_ (
    .A(_03315_),
    .B(_03322_),
    .Y(_03323_)
  );
  AND _11496_ (
    .A(_03308_),
    .B(_03323_),
    .Y(_03324_)
  );
  NAND _11497_ (
    .A(\memory[25][4] ),
    .B(_01469_),
    .Y(_03325_)
  );
  NAND _11498_ (
    .A(\memory[31][4] ),
    .B(_01462_),
    .Y(_03326_)
  );
  AND _11499_ (
    .A(_03325_),
    .B(_03326_),
    .Y(_03327_)
  );
  NAND _11500_ (
    .A(\memory[3][4] ),
    .B(_01449_),
    .Y(_03328_)
  );
  NAND _11501_ (
    .A(\memory[4][4] ),
    .B(_01570_),
    .Y(_03329_)
  );
  AND _11502_ (
    .A(_03328_),
    .B(_03329_),
    .Y(_03330_)
  );
  AND _11503_ (
    .A(_03327_),
    .B(_03330_),
    .Y(_03331_)
  );
  NAND _11504_ (
    .A(\memory[13][4] ),
    .B(_01578_),
    .Y(_03332_)
  );
  NAND _11505_ (
    .A(\memory[16][4] ),
    .B(_01520_),
    .Y(_03333_)
  );
  AND _11506_ (
    .A(_03332_),
    .B(_03333_),
    .Y(_03334_)
  );
  NAND _11507_ (
    .A(\memory[9][4] ),
    .B(_01517_),
    .Y(_03335_)
  );
  NAND _11508_ (
    .A(\memory[5][4] ),
    .B(_01453_),
    .Y(_03336_)
  );
  AND _11509_ (
    .A(_03335_),
    .B(_03336_),
    .Y(_03337_)
  );
  AND _11510_ (
    .A(_03334_),
    .B(_03337_),
    .Y(_03338_)
  );
  AND _11511_ (
    .A(_03331_),
    .B(_03338_),
    .Y(_03339_)
  );
  NAND _11512_ (
    .A(\memory[2][4] ),
    .B(_01504_),
    .Y(_03340_)
  );
  NAND _11513_ (
    .A(\memory[8][4] ),
    .B(_01585_),
    .Y(_03341_)
  );
  AND _11514_ (
    .A(_03340_),
    .B(_03341_),
    .Y(_03342_)
  );
  NAND _11515_ (
    .A(\memory[20][4] ),
    .B(_01479_),
    .Y(_03343_)
  );
  NAND _11516_ (
    .A(\memory[15][4] ),
    .B(_01458_),
    .Y(_03344_)
  );
  AND _11517_ (
    .A(_03343_),
    .B(_03344_),
    .Y(_03345_)
  );
  AND _11518_ (
    .A(_03342_),
    .B(_03345_),
    .Y(_03346_)
  );
  NAND _11519_ (
    .A(\memory[26][4] ),
    .B(_01546_),
    .Y(_03347_)
  );
  NAND _11520_ (
    .A(\memory[27][4] ),
    .B(_01550_),
    .Y(_03348_)
  );
  AND _11521_ (
    .A(_03347_),
    .B(_03348_),
    .Y(_03349_)
  );
  NAND _11522_ (
    .A(\memory[24][4] ),
    .B(_01474_),
    .Y(_03350_)
  );
  NAND _11523_ (
    .A(\memory[6][4] ),
    .B(_01513_),
    .Y(_03351_)
  );
  AND _11524_ (
    .A(_03350_),
    .B(_03351_),
    .Y(_03352_)
  );
  AND _11525_ (
    .A(_03349_),
    .B(_03352_),
    .Y(_03353_)
  );
  AND _11526_ (
    .A(_03346_),
    .B(_03353_),
    .Y(_03354_)
  );
  AND _11527_ (
    .A(_03339_),
    .B(_03354_),
    .Y(_03355_)
  );
  NAND _11528_ (
    .A(_03324_),
    .B(_03355_),
    .Y(_03356_)
  );
  AND _11529_ (
    .A(MemRead_i),
    .B(_03356_),
    .Y(\data_o[28] )
  );
  NAND _11530_ (
    .A(\memory[15][5] ),
    .B(_01458_),
    .Y(_03357_)
  );
  NAND _11531_ (
    .A(\memory[9][5] ),
    .B(_01517_),
    .Y(_03358_)
  );
  AND _11532_ (
    .A(_03357_),
    .B(_03358_),
    .Y(_03359_)
  );
  NAND _11533_ (
    .A(\memory[7][5] ),
    .B(_01530_),
    .Y(_03360_)
  );
  NAND _11534_ (
    .A(\memory[5][5] ),
    .B(_01453_),
    .Y(_03361_)
  );
  AND _11535_ (
    .A(_03360_),
    .B(_03361_),
    .Y(_03362_)
  );
  AND _11536_ (
    .A(_03359_),
    .B(_03362_),
    .Y(_03363_)
  );
  NAND _11537_ (
    .A(\memory[1][5] ),
    .B(_01491_),
    .Y(_03364_)
  );
  NAND _11538_ (
    .A(\memory[8][5] ),
    .B(_01585_),
    .Y(_03365_)
  );
  AND _11539_ (
    .A(_03364_),
    .B(_03365_),
    .Y(_03366_)
  );
  NAND _11540_ (
    .A(\memory[2][5] ),
    .B(_01504_),
    .Y(_03367_)
  );
  NAND _11541_ (
    .A(\memory[31][5] ),
    .B(_01462_),
    .Y(_03368_)
  );
  AND _11542_ (
    .A(_03367_),
    .B(_03368_),
    .Y(_03369_)
  );
  AND _11543_ (
    .A(_03366_),
    .B(_03369_),
    .Y(_03370_)
  );
  AND _11544_ (
    .A(_03363_),
    .B(_03370_),
    .Y(_03371_)
  );
  NAND _11545_ (
    .A(\memory[23][5] ),
    .B(_01553_),
    .Y(_03372_)
  );
  NAND _11546_ (
    .A(\memory[25][5] ),
    .B(_01469_),
    .Y(_03373_)
  );
  AND _11547_ (
    .A(_03372_),
    .B(_03373_),
    .Y(_03374_)
  );
  NAND _11548_ (
    .A(\memory[16][5] ),
    .B(_01520_),
    .Y(_03375_)
  );
  NAND _11549_ (
    .A(\memory[10][5] ),
    .B(_01538_),
    .Y(_03376_)
  );
  AND _11550_ (
    .A(_03375_),
    .B(_03376_),
    .Y(_03377_)
  );
  AND _11551_ (
    .A(_03374_),
    .B(_03377_),
    .Y(_03378_)
  );
  NAND _11552_ (
    .A(\memory[29][5] ),
    .B(_01484_),
    .Y(_03379_)
  );
  NAND _11553_ (
    .A(\memory[21][5] ),
    .B(_01582_),
    .Y(_03380_)
  );
  AND _11554_ (
    .A(_03379_),
    .B(_03380_),
    .Y(_03381_)
  );
  NAND _11555_ (
    .A(\memory[4][5] ),
    .B(_01570_),
    .Y(_03382_)
  );
  NAND _11556_ (
    .A(\memory[3][5] ),
    .B(_01449_),
    .Y(_03383_)
  );
  AND _11557_ (
    .A(_03382_),
    .B(_03383_),
    .Y(_03384_)
  );
  AND _11558_ (
    .A(_03381_),
    .B(_03384_),
    .Y(_03385_)
  );
  AND _11559_ (
    .A(_03378_),
    .B(_03385_),
    .Y(_03386_)
  );
  AND _11560_ (
    .A(_03371_),
    .B(_03386_),
    .Y(_03387_)
  );
  NAND _11561_ (
    .A(\memory[11][5] ),
    .B(_01527_),
    .Y(_03388_)
  );
  NAND _11562_ (
    .A(\memory[19][5] ),
    .B(_01567_),
    .Y(_03389_)
  );
  AND _11563_ (
    .A(_03388_),
    .B(_03389_),
    .Y(_03390_)
  );
  NAND _11564_ (
    .A(\memory[17][5] ),
    .B(_01543_),
    .Y(_03391_)
  );
  NAND _11565_ (
    .A(\memory[6][5] ),
    .B(_01513_),
    .Y(_03392_)
  );
  AND _11566_ (
    .A(_03391_),
    .B(_03392_),
    .Y(_03393_)
  );
  AND _11567_ (
    .A(_03390_),
    .B(_03393_),
    .Y(_03394_)
  );
  NAND _11568_ (
    .A(\memory[14][5] ),
    .B(_01575_),
    .Y(_03395_)
  );
  NAND _11569_ (
    .A(\memory[26][5] ),
    .B(_01546_),
    .Y(_03396_)
  );
  AND _11570_ (
    .A(_03395_),
    .B(_03396_),
    .Y(_03397_)
  );
  NAND _11571_ (
    .A(\memory[12][5] ),
    .B(_01495_),
    .Y(_03398_)
  );
  NAND _11572_ (
    .A(\memory[13][5] ),
    .B(_01578_),
    .Y(_03399_)
  );
  AND _11573_ (
    .A(_03398_),
    .B(_03399_),
    .Y(_03400_)
  );
  AND _11574_ (
    .A(_03397_),
    .B(_03400_),
    .Y(_03401_)
  );
  AND _11575_ (
    .A(_03394_),
    .B(_03401_),
    .Y(_03402_)
  );
  NAND _11576_ (
    .A(\memory[18][5] ),
    .B(_01501_),
    .Y(_03403_)
  );
  NAND _11577_ (
    .A(\memory[20][5] ),
    .B(_01479_),
    .Y(_03404_)
  );
  AND _11578_ (
    .A(_03403_),
    .B(_03404_),
    .Y(_03405_)
  );
  NAND _11579_ (
    .A(\memory[28][5] ),
    .B(_01559_),
    .Y(_03406_)
  );
  NAND _11580_ (
    .A(\memory[0][5] ),
    .B(_01510_),
    .Y(_03407_)
  );
  AND _11581_ (
    .A(_03406_),
    .B(_03407_),
    .Y(_03408_)
  );
  AND _11582_ (
    .A(_03405_),
    .B(_03408_),
    .Y(_03409_)
  );
  NAND _11583_ (
    .A(\memory[27][5] ),
    .B(_01550_),
    .Y(_03410_)
  );
  NAND _11584_ (
    .A(\memory[30][5] ),
    .B(_01563_),
    .Y(_03411_)
  );
  AND _11585_ (
    .A(_03410_),
    .B(_03411_),
    .Y(_03412_)
  );
  NAND _11586_ (
    .A(\memory[24][5] ),
    .B(_01474_),
    .Y(_03413_)
  );
  NAND _11587_ (
    .A(\memory[22][5] ),
    .B(_01534_),
    .Y(_03414_)
  );
  AND _11588_ (
    .A(_03413_),
    .B(_03414_),
    .Y(_03415_)
  );
  AND _11589_ (
    .A(_03412_),
    .B(_03415_),
    .Y(_03416_)
  );
  AND _11590_ (
    .A(_03409_),
    .B(_03416_),
    .Y(_03417_)
  );
  AND _11591_ (
    .A(_03402_),
    .B(_03417_),
    .Y(_03418_)
  );
  NAND _11592_ (
    .A(_03387_),
    .B(_03418_),
    .Y(_03419_)
  );
  AND _11593_ (
    .A(MemRead_i),
    .B(_03419_),
    .Y(\data_o[29] )
  );
  NAND _11594_ (
    .A(\memory[12][6] ),
    .B(_01495_),
    .Y(_03420_)
  );
  NAND _11595_ (
    .A(\memory[2][6] ),
    .B(_01504_),
    .Y(_03421_)
  );
  AND _11596_ (
    .A(_03420_),
    .B(_03421_),
    .Y(_03422_)
  );
  NAND _11597_ (
    .A(\memory[4][6] ),
    .B(_01570_),
    .Y(_03423_)
  );
  NAND _11598_ (
    .A(\memory[8][6] ),
    .B(_01585_),
    .Y(_03424_)
  );
  AND _11599_ (
    .A(_03423_),
    .B(_03424_),
    .Y(_03425_)
  );
  AND _11600_ (
    .A(_03422_),
    .B(_03425_),
    .Y(_03426_)
  );
  NAND _11601_ (
    .A(\memory[16][6] ),
    .B(_01520_),
    .Y(_03427_)
  );
  NAND _11602_ (
    .A(\memory[15][6] ),
    .B(_01458_),
    .Y(_03428_)
  );
  AND _11603_ (
    .A(_03427_),
    .B(_03428_),
    .Y(_03429_)
  );
  NAND _11604_ (
    .A(\memory[25][6] ),
    .B(_01469_),
    .Y(_03430_)
  );
  NAND _11605_ (
    .A(\memory[14][6] ),
    .B(_01575_),
    .Y(_03431_)
  );
  AND _11606_ (
    .A(_03430_),
    .B(_03431_),
    .Y(_03432_)
  );
  AND _11607_ (
    .A(_03429_),
    .B(_03432_),
    .Y(_03433_)
  );
  AND _11608_ (
    .A(_03426_),
    .B(_03433_),
    .Y(_03434_)
  );
  NAND _11609_ (
    .A(\memory[10][6] ),
    .B(_01538_),
    .Y(_03435_)
  );
  NAND _11610_ (
    .A(\memory[3][6] ),
    .B(_01449_),
    .Y(_03436_)
  );
  AND _11611_ (
    .A(_03435_),
    .B(_03436_),
    .Y(_03437_)
  );
  NAND _11612_ (
    .A(\memory[5][6] ),
    .B(_01453_),
    .Y(_03438_)
  );
  NAND _11613_ (
    .A(\memory[29][6] ),
    .B(_01484_),
    .Y(_03439_)
  );
  AND _11614_ (
    .A(_03438_),
    .B(_03439_),
    .Y(_03440_)
  );
  AND _11615_ (
    .A(_03437_),
    .B(_03440_),
    .Y(_03441_)
  );
  NAND _11616_ (
    .A(\memory[13][6] ),
    .B(_01578_),
    .Y(_03442_)
  );
  NAND _11617_ (
    .A(\memory[30][6] ),
    .B(_01563_),
    .Y(_03443_)
  );
  AND _11618_ (
    .A(_03442_),
    .B(_03443_),
    .Y(_03444_)
  );
  NAND _11619_ (
    .A(\memory[18][6] ),
    .B(_01501_),
    .Y(_03445_)
  );
  NAND _11620_ (
    .A(\memory[22][6] ),
    .B(_01534_),
    .Y(_03446_)
  );
  AND _11621_ (
    .A(_03445_),
    .B(_03446_),
    .Y(_03447_)
  );
  AND _11622_ (
    .A(_03444_),
    .B(_03447_),
    .Y(_03448_)
  );
  AND _11623_ (
    .A(_03441_),
    .B(_03448_),
    .Y(_03449_)
  );
  AND _11624_ (
    .A(_03434_),
    .B(_03449_),
    .Y(_03450_)
  );
  NAND _11625_ (
    .A(\memory[9][6] ),
    .B(_01517_),
    .Y(_03451_)
  );
  NAND _11626_ (
    .A(\memory[1][6] ),
    .B(_01491_),
    .Y(_03452_)
  );
  AND _11627_ (
    .A(_03451_),
    .B(_03452_),
    .Y(_03453_)
  );
  NAND _11628_ (
    .A(\memory[21][6] ),
    .B(_01582_),
    .Y(_03454_)
  );
  NAND _11629_ (
    .A(\memory[7][6] ),
    .B(_01530_),
    .Y(_03455_)
  );
  AND _11630_ (
    .A(_03454_),
    .B(_03455_),
    .Y(_03456_)
  );
  AND _11631_ (
    .A(_03453_),
    .B(_03456_),
    .Y(_03457_)
  );
  NAND _11632_ (
    .A(\memory[23][6] ),
    .B(_01553_),
    .Y(_03458_)
  );
  NAND _11633_ (
    .A(\memory[6][6] ),
    .B(_01513_),
    .Y(_03459_)
  );
  AND _11634_ (
    .A(_03458_),
    .B(_03459_),
    .Y(_03460_)
  );
  NAND _11635_ (
    .A(\memory[24][6] ),
    .B(_01474_),
    .Y(_03461_)
  );
  NAND _11636_ (
    .A(\memory[19][6] ),
    .B(_01567_),
    .Y(_03462_)
  );
  AND _11637_ (
    .A(_03461_),
    .B(_03462_),
    .Y(_03463_)
  );
  AND _11638_ (
    .A(_03460_),
    .B(_03463_),
    .Y(_03464_)
  );
  AND _11639_ (
    .A(_03457_),
    .B(_03464_),
    .Y(_03465_)
  );
  NAND _11640_ (
    .A(\memory[31][6] ),
    .B(_01462_),
    .Y(_03466_)
  );
  NAND _11641_ (
    .A(\memory[28][6] ),
    .B(_01559_),
    .Y(_03467_)
  );
  AND _11642_ (
    .A(_03466_),
    .B(_03467_),
    .Y(_03468_)
  );
  NAND _11643_ (
    .A(\memory[17][6] ),
    .B(_01543_),
    .Y(_03469_)
  );
  NAND _11644_ (
    .A(\memory[11][6] ),
    .B(_01527_),
    .Y(_03470_)
  );
  AND _11645_ (
    .A(_03469_),
    .B(_03470_),
    .Y(_03471_)
  );
  AND _11646_ (
    .A(_03468_),
    .B(_03471_),
    .Y(_03472_)
  );
  NAND _11647_ (
    .A(\memory[27][6] ),
    .B(_01550_),
    .Y(_03473_)
  );
  NAND _11648_ (
    .A(\memory[0][6] ),
    .B(_01510_),
    .Y(_03474_)
  );
  AND _11649_ (
    .A(_03473_),
    .B(_03474_),
    .Y(_03475_)
  );
  NAND _11650_ (
    .A(\memory[20][6] ),
    .B(_01479_),
    .Y(_03476_)
  );
  NAND _11651_ (
    .A(\memory[26][6] ),
    .B(_01546_),
    .Y(_03477_)
  );
  AND _11652_ (
    .A(_03476_),
    .B(_03477_),
    .Y(_03478_)
  );
  AND _11653_ (
    .A(_03475_),
    .B(_03478_),
    .Y(_03479_)
  );
  AND _11654_ (
    .A(_03472_),
    .B(_03479_),
    .Y(_03480_)
  );
  AND _11655_ (
    .A(_03465_),
    .B(_03480_),
    .Y(_03481_)
  );
  NAND _11656_ (
    .A(_03450_),
    .B(_03481_),
    .Y(_03482_)
  );
  AND _11657_ (
    .A(MemRead_i),
    .B(_03482_),
    .Y(\data_o[30] )
  );
  NAND _11658_ (
    .A(\memory[27][7] ),
    .B(_01550_),
    .Y(_03483_)
  );
  NAND _11659_ (
    .A(\memory[0][7] ),
    .B(_01510_),
    .Y(_03484_)
  );
  AND _11660_ (
    .A(_03483_),
    .B(_03484_),
    .Y(_03485_)
  );
  NAND _11661_ (
    .A(\memory[31][7] ),
    .B(_01462_),
    .Y(_03486_)
  );
  NAND _11662_ (
    .A(\memory[18][7] ),
    .B(_01501_),
    .Y(_03487_)
  );
  AND _11663_ (
    .A(_03486_),
    .B(_03487_),
    .Y(_03488_)
  );
  AND _11664_ (
    .A(_03485_),
    .B(_03488_),
    .Y(_03489_)
  );
  NAND _11665_ (
    .A(\memory[28][7] ),
    .B(_01559_),
    .Y(_03490_)
  );
  NAND _11666_ (
    .A(\memory[25][7] ),
    .B(_01469_),
    .Y(_03491_)
  );
  AND _11667_ (
    .A(_03490_),
    .B(_03491_),
    .Y(_03492_)
  );
  NAND _11668_ (
    .A(\memory[19][7] ),
    .B(_01567_),
    .Y(_03493_)
  );
  NAND _11669_ (
    .A(\memory[3][7] ),
    .B(_01449_),
    .Y(_03494_)
  );
  AND _11670_ (
    .A(_03493_),
    .B(_03494_),
    .Y(_03495_)
  );
  AND _11671_ (
    .A(_03492_),
    .B(_03495_),
    .Y(_03496_)
  );
  AND _11672_ (
    .A(_03489_),
    .B(_03496_),
    .Y(_03497_)
  );
  NAND _11673_ (
    .A(\memory[9][7] ),
    .B(_01517_),
    .Y(_03498_)
  );
  NAND _11674_ (
    .A(\memory[4][7] ),
    .B(_01570_),
    .Y(_03499_)
  );
  AND _11675_ (
    .A(_03498_),
    .B(_03499_),
    .Y(_03500_)
  );
  NAND _11676_ (
    .A(\memory[30][7] ),
    .B(_01563_),
    .Y(_03501_)
  );
  NAND _11677_ (
    .A(\memory[7][7] ),
    .B(_01530_),
    .Y(_03502_)
  );
  AND _11678_ (
    .A(_03501_),
    .B(_03502_),
    .Y(_03503_)
  );
  AND _11679_ (
    .A(_03500_),
    .B(_03503_),
    .Y(_03504_)
  );
  NAND _11680_ (
    .A(\memory[29][7] ),
    .B(_01484_),
    .Y(_03505_)
  );
  NAND _11681_ (
    .A(\memory[1][7] ),
    .B(_01491_),
    .Y(_03506_)
  );
  AND _11682_ (
    .A(_03505_),
    .B(_03506_),
    .Y(_03507_)
  );
  NAND _11683_ (
    .A(\memory[13][7] ),
    .B(_01578_),
    .Y(_03508_)
  );
  NAND _11684_ (
    .A(\memory[20][7] ),
    .B(_01479_),
    .Y(_03509_)
  );
  AND _11685_ (
    .A(_03508_),
    .B(_03509_),
    .Y(_03510_)
  );
  AND _11686_ (
    .A(_03507_),
    .B(_03510_),
    .Y(_03511_)
  );
  AND _11687_ (
    .A(_03504_),
    .B(_03511_),
    .Y(_03512_)
  );
  AND _11688_ (
    .A(_03497_),
    .B(_03512_),
    .Y(_03513_)
  );
  NAND _11689_ (
    .A(\memory[2][7] ),
    .B(_01504_),
    .Y(_03514_)
  );
  NAND _11690_ (
    .A(\memory[12][7] ),
    .B(_01495_),
    .Y(_03515_)
  );
  AND _11691_ (
    .A(_03514_),
    .B(_03515_),
    .Y(_03516_)
  );
  NAND _11692_ (
    .A(\memory[11][7] ),
    .B(_01527_),
    .Y(_03517_)
  );
  NAND _11693_ (
    .A(\memory[23][7] ),
    .B(_01553_),
    .Y(_03518_)
  );
  AND _11694_ (
    .A(_03517_),
    .B(_03518_),
    .Y(_03519_)
  );
  AND _11695_ (
    .A(_03516_),
    .B(_03519_),
    .Y(_03520_)
  );
  NAND _11696_ (
    .A(\memory[6][7] ),
    .B(_01513_),
    .Y(_03521_)
  );
  NAND _11697_ (
    .A(\memory[5][7] ),
    .B(_01453_),
    .Y(_03522_)
  );
  AND _11698_ (
    .A(_03521_),
    .B(_03522_),
    .Y(_03523_)
  );
  NAND _11699_ (
    .A(\memory[16][7] ),
    .B(_01520_),
    .Y(_03524_)
  );
  NAND _11700_ (
    .A(\memory[22][7] ),
    .B(_01534_),
    .Y(_03525_)
  );
  AND _11701_ (
    .A(_03524_),
    .B(_03525_),
    .Y(_03526_)
  );
  AND _11702_ (
    .A(_03523_),
    .B(_03526_),
    .Y(_03527_)
  );
  AND _11703_ (
    .A(_03520_),
    .B(_03527_),
    .Y(_03528_)
  );
  NAND _11704_ (
    .A(\memory[21][7] ),
    .B(_01582_),
    .Y(_03529_)
  );
  NAND _11705_ (
    .A(\memory[24][7] ),
    .B(_01474_),
    .Y(_03530_)
  );
  AND _11706_ (
    .A(_03529_),
    .B(_03530_),
    .Y(_03531_)
  );
  NAND _11707_ (
    .A(\memory[17][7] ),
    .B(_01543_),
    .Y(_03532_)
  );
  NAND _11708_ (
    .A(\memory[26][7] ),
    .B(_01546_),
    .Y(_03533_)
  );
  AND _11709_ (
    .A(_03532_),
    .B(_03533_),
    .Y(_03534_)
  );
  AND _11710_ (
    .A(_03531_),
    .B(_03534_),
    .Y(_03535_)
  );
  NAND _11711_ (
    .A(\memory[8][7] ),
    .B(_01585_),
    .Y(_03536_)
  );
  NAND _11712_ (
    .A(\memory[10][7] ),
    .B(_01538_),
    .Y(_03537_)
  );
  AND _11713_ (
    .A(_03536_),
    .B(_03537_),
    .Y(_03538_)
  );
  NAND _11714_ (
    .A(\memory[14][7] ),
    .B(_01575_),
    .Y(_03539_)
  );
  NAND _11715_ (
    .A(\memory[15][7] ),
    .B(_01458_),
    .Y(_03540_)
  );
  AND _11716_ (
    .A(_03539_),
    .B(_03540_),
    .Y(_03541_)
  );
  AND _11717_ (
    .A(_03538_),
    .B(_03541_),
    .Y(_03542_)
  );
  AND _11718_ (
    .A(_03535_),
    .B(_03542_),
    .Y(_03543_)
  );
  AND _11719_ (
    .A(_03528_),
    .B(_03543_),
    .Y(_03544_)
  );
  NAND _11720_ (
    .A(_03513_),
    .B(_03544_),
    .Y(_03545_)
  );
  AND _11721_ (
    .A(MemRead_i),
    .B(_03545_),
    .Y(\data_o[31] )
  );
  NAND _11722_ (
    .A(\memory[31][0] ),
    .B(_05361_),
    .Y(_03546_)
  );
  OR _11723_ (
    .A(\memory[31][0] ),
    .B(_01462_),
    .Y(_03547_)
  );
  OR _11724_ (
    .A(\data_i[24] ),
    .B(_01463_),
    .Y(_03548_)
  );
  NAND _11725_ (
    .A(_03547_),
    .B(_03548_),
    .Y(_03549_)
  );
  NAND _11726_ (
    .A(_01511_),
    .B(_03549_),
    .Y(_03550_)
  );
  OR _11727_ (
    .A(\data_i[16] ),
    .B(_01511_),
    .Y(_03551_)
  );
  AND _11728_ (
    .A(_03550_),
    .B(_03551_),
    .Y(_03552_)
  );
  NAND _11729_ (
    .A(\data_i[8] ),
    .B(_01491_),
    .Y(_03553_)
  );
  AND _11730_ (
    .A(_01505_),
    .B(_03553_),
    .Y(_03554_)
  );
  NAND _11731_ (
    .A(_01492_),
    .B(_03552_),
    .Y(_03555_)
  );
  NAND _11732_ (
    .A(_03554_),
    .B(_03555_),
    .Y(_03556_)
  );
  OR _11733_ (
    .A(\data_i[0] ),
    .B(_01505_),
    .Y(_03557_)
  );
  AND _11734_ (
    .A(MemWrite_i),
    .B(_03557_),
    .Y(_03558_)
  );
  NAND _11735_ (
    .A(_03556_),
    .B(_03558_),
    .Y(_03559_)
  );
  NAND _11736_ (
    .A(_03546_),
    .B(_03559_),
    .Y(_00192_)
  );
  NAND _11737_ (
    .A(\memory[31][1] ),
    .B(_05361_),
    .Y(_03560_)
  );
  OR _11738_ (
    .A(\memory[31][1] ),
    .B(_01462_),
    .Y(_03561_)
  );
  OR _11739_ (
    .A(\data_i[25] ),
    .B(_01463_),
    .Y(_03562_)
  );
  NAND _11740_ (
    .A(_03561_),
    .B(_03562_),
    .Y(_03563_)
  );
  NAND _11741_ (
    .A(_01511_),
    .B(_03563_),
    .Y(_03564_)
  );
  OR _11742_ (
    .A(\data_i[17] ),
    .B(_01511_),
    .Y(_03565_)
  );
  AND _11743_ (
    .A(_03564_),
    .B(_03565_),
    .Y(_03566_)
  );
  NAND _11744_ (
    .A(\data_i[9] ),
    .B(_01491_),
    .Y(_03567_)
  );
  AND _11745_ (
    .A(_01505_),
    .B(_03567_),
    .Y(_03568_)
  );
  NAND _11746_ (
    .A(_01492_),
    .B(_03566_),
    .Y(_03569_)
  );
  NAND _11747_ (
    .A(_03568_),
    .B(_03569_),
    .Y(_03570_)
  );
  OR _11748_ (
    .A(\data_i[1] ),
    .B(_01505_),
    .Y(_03571_)
  );
  AND _11749_ (
    .A(MemWrite_i),
    .B(_03571_),
    .Y(_03572_)
  );
  NAND _11750_ (
    .A(_03570_),
    .B(_03572_),
    .Y(_03573_)
  );
  NAND _11751_ (
    .A(_03560_),
    .B(_03573_),
    .Y(_00193_)
  );
  NAND _11752_ (
    .A(\memory[31][2] ),
    .B(_05361_),
    .Y(_03574_)
  );
  OR _11753_ (
    .A(\memory[31][2] ),
    .B(_01462_),
    .Y(_03575_)
  );
  OR _11754_ (
    .A(\data_i[26] ),
    .B(_01463_),
    .Y(_03576_)
  );
  NAND _11755_ (
    .A(_03575_),
    .B(_03576_),
    .Y(_03577_)
  );
  NAND _11756_ (
    .A(_01511_),
    .B(_03577_),
    .Y(_03578_)
  );
  OR _11757_ (
    .A(\data_i[18] ),
    .B(_01511_),
    .Y(_03579_)
  );
  AND _11758_ (
    .A(_03578_),
    .B(_03579_),
    .Y(_03580_)
  );
  NAND _11759_ (
    .A(\data_i[10] ),
    .B(_01491_),
    .Y(_03581_)
  );
  AND _11760_ (
    .A(_01505_),
    .B(_03581_),
    .Y(_03582_)
  );
  NAND _11761_ (
    .A(_01492_),
    .B(_03580_),
    .Y(_03583_)
  );
  NAND _11762_ (
    .A(_03582_),
    .B(_03583_),
    .Y(_03584_)
  );
  OR _11763_ (
    .A(\data_i[2] ),
    .B(_01505_),
    .Y(_03585_)
  );
  AND _11764_ (
    .A(MemWrite_i),
    .B(_03585_),
    .Y(_03586_)
  );
  NAND _11765_ (
    .A(_03584_),
    .B(_03586_),
    .Y(_03587_)
  );
  NAND _11766_ (
    .A(_03574_),
    .B(_03587_),
    .Y(_00194_)
  );
  NAND _11767_ (
    .A(\memory[31][3] ),
    .B(_05361_),
    .Y(_03588_)
  );
  OR _11768_ (
    .A(\memory[31][3] ),
    .B(_01462_),
    .Y(_03589_)
  );
  OR _11769_ (
    .A(\data_i[27] ),
    .B(_01463_),
    .Y(_03590_)
  );
  NAND _11770_ (
    .A(_03589_),
    .B(_03590_),
    .Y(_03591_)
  );
  NAND _11771_ (
    .A(_01511_),
    .B(_03591_),
    .Y(_03592_)
  );
  OR _11772_ (
    .A(\data_i[19] ),
    .B(_01511_),
    .Y(_03593_)
  );
  AND _11773_ (
    .A(_03592_),
    .B(_03593_),
    .Y(_03594_)
  );
  NAND _11774_ (
    .A(\data_i[11] ),
    .B(_01491_),
    .Y(_03595_)
  );
  AND _11775_ (
    .A(_01505_),
    .B(_03595_),
    .Y(_03596_)
  );
  NAND _11776_ (
    .A(_01492_),
    .B(_03594_),
    .Y(_03597_)
  );
  NAND _11777_ (
    .A(_03596_),
    .B(_03597_),
    .Y(_03598_)
  );
  OR _11778_ (
    .A(\data_i[3] ),
    .B(_01505_),
    .Y(_03599_)
  );
  AND _11779_ (
    .A(MemWrite_i),
    .B(_03599_),
    .Y(_03600_)
  );
  NAND _11780_ (
    .A(_03598_),
    .B(_03600_),
    .Y(_03601_)
  );
  NAND _11781_ (
    .A(_03588_),
    .B(_03601_),
    .Y(_00195_)
  );
  NAND _11782_ (
    .A(\memory[31][4] ),
    .B(_05361_),
    .Y(_03602_)
  );
  OR _11783_ (
    .A(\memory[31][4] ),
    .B(_01462_),
    .Y(_03603_)
  );
  OR _11784_ (
    .A(\data_i[28] ),
    .B(_01463_),
    .Y(_03604_)
  );
  NAND _11785_ (
    .A(_03603_),
    .B(_03604_),
    .Y(_03605_)
  );
  NAND _11786_ (
    .A(_01511_),
    .B(_03605_),
    .Y(_03606_)
  );
  OR _11787_ (
    .A(\data_i[20] ),
    .B(_01511_),
    .Y(_03607_)
  );
  AND _11788_ (
    .A(_03606_),
    .B(_03607_),
    .Y(_03608_)
  );
  NAND _11789_ (
    .A(\data_i[12] ),
    .B(_01491_),
    .Y(_03609_)
  );
  AND _11790_ (
    .A(_01505_),
    .B(_03609_),
    .Y(_03610_)
  );
  NAND _11791_ (
    .A(_01492_),
    .B(_03608_),
    .Y(_03611_)
  );
  NAND _11792_ (
    .A(_03610_),
    .B(_03611_),
    .Y(_03612_)
  );
  OR _11793_ (
    .A(\data_i[4] ),
    .B(_01505_),
    .Y(_03613_)
  );
  AND _11794_ (
    .A(MemWrite_i),
    .B(_03613_),
    .Y(_03614_)
  );
  NAND _11795_ (
    .A(_03612_),
    .B(_03614_),
    .Y(_03615_)
  );
  NAND _11796_ (
    .A(_03602_),
    .B(_03615_),
    .Y(_00196_)
  );
  NAND _11797_ (
    .A(\memory[31][5] ),
    .B(_05361_),
    .Y(_03616_)
  );
  OR _11798_ (
    .A(\memory[31][5] ),
    .B(_01462_),
    .Y(_03617_)
  );
  OR _11799_ (
    .A(\data_i[29] ),
    .B(_01463_),
    .Y(_03618_)
  );
  NAND _11800_ (
    .A(_03617_),
    .B(_03618_),
    .Y(_03619_)
  );
  NAND _11801_ (
    .A(_01511_),
    .B(_03619_),
    .Y(_03620_)
  );
  OR _11802_ (
    .A(\data_i[21] ),
    .B(_01511_),
    .Y(_03621_)
  );
  AND _11803_ (
    .A(_03620_),
    .B(_03621_),
    .Y(_03622_)
  );
  NAND _11804_ (
    .A(\data_i[13] ),
    .B(_01491_),
    .Y(_03623_)
  );
  AND _11805_ (
    .A(_01505_),
    .B(_03623_),
    .Y(_03624_)
  );
  NAND _11806_ (
    .A(_01492_),
    .B(_03622_),
    .Y(_03625_)
  );
  NAND _11807_ (
    .A(_03624_),
    .B(_03625_),
    .Y(_03626_)
  );
  OR _11808_ (
    .A(\data_i[5] ),
    .B(_01505_),
    .Y(_03627_)
  );
  AND _11809_ (
    .A(MemWrite_i),
    .B(_03627_),
    .Y(_03628_)
  );
  NAND _11810_ (
    .A(_03626_),
    .B(_03628_),
    .Y(_03629_)
  );
  NAND _11811_ (
    .A(_03616_),
    .B(_03629_),
    .Y(_00197_)
  );
  NAND _11812_ (
    .A(\memory[31][6] ),
    .B(_05361_),
    .Y(_03630_)
  );
  OR _11813_ (
    .A(\memory[31][6] ),
    .B(_01462_),
    .Y(_03631_)
  );
  OR _11814_ (
    .A(\data_i[30] ),
    .B(_01463_),
    .Y(_03632_)
  );
  NAND _11815_ (
    .A(_03631_),
    .B(_03632_),
    .Y(_03633_)
  );
  NAND _11816_ (
    .A(_01511_),
    .B(_03633_),
    .Y(_03634_)
  );
  OR _11817_ (
    .A(\data_i[22] ),
    .B(_01511_),
    .Y(_03635_)
  );
  AND _11818_ (
    .A(_03634_),
    .B(_03635_),
    .Y(_03636_)
  );
  NAND _11819_ (
    .A(\data_i[14] ),
    .B(_01491_),
    .Y(_03637_)
  );
  AND _11820_ (
    .A(_01505_),
    .B(_03637_),
    .Y(_03638_)
  );
  NAND _11821_ (
    .A(_01492_),
    .B(_03636_),
    .Y(_03639_)
  );
  NAND _11822_ (
    .A(_03638_),
    .B(_03639_),
    .Y(_03640_)
  );
  OR _11823_ (
    .A(\data_i[6] ),
    .B(_01505_),
    .Y(_03641_)
  );
  AND _11824_ (
    .A(MemWrite_i),
    .B(_03641_),
    .Y(_03642_)
  );
  NAND _11825_ (
    .A(_03640_),
    .B(_03642_),
    .Y(_03643_)
  );
  NAND _11826_ (
    .A(_03630_),
    .B(_03643_),
    .Y(_00198_)
  );
  NAND _11827_ (
    .A(\memory[31][7] ),
    .B(_05361_),
    .Y(_03644_)
  );
  OR _11828_ (
    .A(\memory[31][7] ),
    .B(_01462_),
    .Y(_03645_)
  );
  OR _11829_ (
    .A(\data_i[31] ),
    .B(_01463_),
    .Y(_03646_)
  );
  NAND _11830_ (
    .A(_03645_),
    .B(_03646_),
    .Y(_03647_)
  );
  NAND _11831_ (
    .A(_01511_),
    .B(_03647_),
    .Y(_03648_)
  );
  OR _11832_ (
    .A(\data_i[23] ),
    .B(_01511_),
    .Y(_03649_)
  );
  AND _11833_ (
    .A(_03648_),
    .B(_03649_),
    .Y(_03650_)
  );
  NAND _11834_ (
    .A(\data_i[15] ),
    .B(_01491_),
    .Y(_03651_)
  );
  AND _11835_ (
    .A(_01505_),
    .B(_03651_),
    .Y(_03652_)
  );
  NAND _11836_ (
    .A(_01492_),
    .B(_03650_),
    .Y(_03653_)
  );
  NAND _11837_ (
    .A(_03652_),
    .B(_03653_),
    .Y(_03654_)
  );
  OR _11838_ (
    .A(\data_i[7] ),
    .B(_01505_),
    .Y(_03655_)
  );
  AND _11839_ (
    .A(MemWrite_i),
    .B(_03655_),
    .Y(_03656_)
  );
  NAND _11840_ (
    .A(_03654_),
    .B(_03656_),
    .Y(_03657_)
  );
  NAND _11841_ (
    .A(_03644_),
    .B(_03657_),
    .Y(_00199_)
  );
  NAND _11842_ (
    .A(\memory[30][0] ),
    .B(_05361_),
    .Y(_03658_)
  );
  OR _11843_ (
    .A(\memory[30][0] ),
    .B(_01563_),
    .Y(_03659_)
  );
  OR _11844_ (
    .A(\data_i[24] ),
    .B(_01564_),
    .Y(_03660_)
  );
  NAND _11845_ (
    .A(_03659_),
    .B(_03660_),
    .Y(_03661_)
  );
  NAND _11846_ (
    .A(_01463_),
    .B(_03661_),
    .Y(_03662_)
  );
  OR _11847_ (
    .A(\data_i[16] ),
    .B(_01463_),
    .Y(_03663_)
  );
  AND _11848_ (
    .A(_03662_),
    .B(_03663_),
    .Y(_03664_)
  );
  NAND _11849_ (
    .A(\data_i[8] ),
    .B(_01510_),
    .Y(_03665_)
  );
  AND _11850_ (
    .A(_01492_),
    .B(_03665_),
    .Y(_03666_)
  );
  NAND _11851_ (
    .A(_01511_),
    .B(_03664_),
    .Y(_03667_)
  );
  NAND _11852_ (
    .A(_03666_),
    .B(_03667_),
    .Y(_03668_)
  );
  OR _11853_ (
    .A(\data_i[0] ),
    .B(_01492_),
    .Y(_03669_)
  );
  AND _11854_ (
    .A(MemWrite_i),
    .B(_03669_),
    .Y(_03670_)
  );
  NAND _11855_ (
    .A(_03668_),
    .B(_03670_),
    .Y(_03671_)
  );
  NAND _11856_ (
    .A(_03658_),
    .B(_03671_),
    .Y(_00184_)
  );
  NAND _11857_ (
    .A(\memory[30][1] ),
    .B(_05361_),
    .Y(_03672_)
  );
  OR _11858_ (
    .A(\memory[30][1] ),
    .B(_01563_),
    .Y(_03673_)
  );
  OR _11859_ (
    .A(\data_i[25] ),
    .B(_01564_),
    .Y(_03674_)
  );
  NAND _11860_ (
    .A(_03673_),
    .B(_03674_),
    .Y(_03675_)
  );
  NAND _11861_ (
    .A(_01463_),
    .B(_03675_),
    .Y(_03676_)
  );
  OR _11862_ (
    .A(\data_i[17] ),
    .B(_01463_),
    .Y(_03677_)
  );
  AND _11863_ (
    .A(_03676_),
    .B(_03677_),
    .Y(_03678_)
  );
  NAND _11864_ (
    .A(\data_i[9] ),
    .B(_01510_),
    .Y(_03679_)
  );
  AND _11865_ (
    .A(_01492_),
    .B(_03679_),
    .Y(_03680_)
  );
  NAND _11866_ (
    .A(_01511_),
    .B(_03678_),
    .Y(_03681_)
  );
  NAND _11867_ (
    .A(_03680_),
    .B(_03681_),
    .Y(_03682_)
  );
  OR _11868_ (
    .A(\data_i[1] ),
    .B(_01492_),
    .Y(_03683_)
  );
  AND _11869_ (
    .A(MemWrite_i),
    .B(_03683_),
    .Y(_03684_)
  );
  NAND _11870_ (
    .A(_03682_),
    .B(_03684_),
    .Y(_03685_)
  );
  NAND _11871_ (
    .A(_03672_),
    .B(_03685_),
    .Y(_00185_)
  );
  NAND _11872_ (
    .A(\memory[30][2] ),
    .B(_05361_),
    .Y(_03686_)
  );
  OR _11873_ (
    .A(\memory[30][2] ),
    .B(_01563_),
    .Y(_03687_)
  );
  OR _11874_ (
    .A(\data_i[26] ),
    .B(_01564_),
    .Y(_03688_)
  );
  NAND _11875_ (
    .A(_03687_),
    .B(_03688_),
    .Y(_03689_)
  );
  NAND _11876_ (
    .A(_01463_),
    .B(_03689_),
    .Y(_03690_)
  );
  OR _11877_ (
    .A(\data_i[18] ),
    .B(_01463_),
    .Y(_03691_)
  );
  AND _11878_ (
    .A(_03690_),
    .B(_03691_),
    .Y(_03692_)
  );
  NAND _11879_ (
    .A(\data_i[10] ),
    .B(_01510_),
    .Y(_03693_)
  );
  AND _11880_ (
    .A(_01492_),
    .B(_03693_),
    .Y(_03694_)
  );
  NAND _11881_ (
    .A(_01511_),
    .B(_03692_),
    .Y(_03695_)
  );
  NAND _11882_ (
    .A(_03694_),
    .B(_03695_),
    .Y(_03696_)
  );
  OR _11883_ (
    .A(\data_i[2] ),
    .B(_01492_),
    .Y(_03697_)
  );
  AND _11884_ (
    .A(MemWrite_i),
    .B(_03697_),
    .Y(_03698_)
  );
  NAND _11885_ (
    .A(_03696_),
    .B(_03698_),
    .Y(_03699_)
  );
  NAND _11886_ (
    .A(_03686_),
    .B(_03699_),
    .Y(_00186_)
  );
  NAND _11887_ (
    .A(\memory[30][3] ),
    .B(_05361_),
    .Y(_03700_)
  );
  OR _11888_ (
    .A(\memory[30][3] ),
    .B(_01563_),
    .Y(_03701_)
  );
  OR _11889_ (
    .A(\data_i[27] ),
    .B(_01564_),
    .Y(_03702_)
  );
  NAND _11890_ (
    .A(_03701_),
    .B(_03702_),
    .Y(_03703_)
  );
  NAND _11891_ (
    .A(_01463_),
    .B(_03703_),
    .Y(_03704_)
  );
  OR _11892_ (
    .A(\data_i[19] ),
    .B(_01463_),
    .Y(_03705_)
  );
  AND _11893_ (
    .A(_03704_),
    .B(_03705_),
    .Y(_03706_)
  );
  NAND _11894_ (
    .A(\data_i[11] ),
    .B(_01510_),
    .Y(_03707_)
  );
  AND _11895_ (
    .A(_01492_),
    .B(_03707_),
    .Y(_03708_)
  );
  NAND _11896_ (
    .A(_01511_),
    .B(_03706_),
    .Y(_03709_)
  );
  NAND _11897_ (
    .A(_03708_),
    .B(_03709_),
    .Y(_03710_)
  );
  OR _11898_ (
    .A(\data_i[3] ),
    .B(_01492_),
    .Y(_03711_)
  );
  AND _11899_ (
    .A(MemWrite_i),
    .B(_03711_),
    .Y(_03712_)
  );
  NAND _11900_ (
    .A(_03710_),
    .B(_03712_),
    .Y(_03713_)
  );
  NAND _11901_ (
    .A(_03700_),
    .B(_03713_),
    .Y(_00187_)
  );
  NAND _11902_ (
    .A(\memory[30][4] ),
    .B(_05361_),
    .Y(_03714_)
  );
  OR _11903_ (
    .A(\memory[30][4] ),
    .B(_01563_),
    .Y(_03715_)
  );
  OR _11904_ (
    .A(\data_i[28] ),
    .B(_01564_),
    .Y(_03716_)
  );
  NAND _11905_ (
    .A(_03715_),
    .B(_03716_),
    .Y(_03717_)
  );
  NAND _11906_ (
    .A(_01463_),
    .B(_03717_),
    .Y(_03718_)
  );
  OR _11907_ (
    .A(\data_i[20] ),
    .B(_01463_),
    .Y(_03719_)
  );
  AND _11908_ (
    .A(_03718_),
    .B(_03719_),
    .Y(_03720_)
  );
  NAND _11909_ (
    .A(\data_i[12] ),
    .B(_01510_),
    .Y(_03721_)
  );
  AND _11910_ (
    .A(_01492_),
    .B(_03721_),
    .Y(_03722_)
  );
  NAND _11911_ (
    .A(_01511_),
    .B(_03720_),
    .Y(_03723_)
  );
  NAND _11912_ (
    .A(_03722_),
    .B(_03723_),
    .Y(_03724_)
  );
  OR _11913_ (
    .A(\data_i[4] ),
    .B(_01492_),
    .Y(_03725_)
  );
  AND _11914_ (
    .A(MemWrite_i),
    .B(_03725_),
    .Y(_03726_)
  );
  NAND _11915_ (
    .A(_03724_),
    .B(_03726_),
    .Y(_03727_)
  );
  NAND _11916_ (
    .A(_03714_),
    .B(_03727_),
    .Y(_00188_)
  );
  NAND _11917_ (
    .A(\memory[30][5] ),
    .B(_05361_),
    .Y(_03728_)
  );
  OR _11918_ (
    .A(\memory[30][5] ),
    .B(_01563_),
    .Y(_03729_)
  );
  OR _11919_ (
    .A(\data_i[29] ),
    .B(_01564_),
    .Y(_03730_)
  );
  NAND _11920_ (
    .A(_03729_),
    .B(_03730_),
    .Y(_03731_)
  );
  NAND _11921_ (
    .A(_01463_),
    .B(_03731_),
    .Y(_03732_)
  );
  OR _11922_ (
    .A(\data_i[21] ),
    .B(_01463_),
    .Y(_03733_)
  );
  AND _11923_ (
    .A(_03732_),
    .B(_03733_),
    .Y(_03734_)
  );
  NAND _11924_ (
    .A(\data_i[13] ),
    .B(_01510_),
    .Y(_03735_)
  );
  AND _11925_ (
    .A(_01492_),
    .B(_03735_),
    .Y(_03736_)
  );
  NAND _11926_ (
    .A(_01511_),
    .B(_03734_),
    .Y(_03737_)
  );
  NAND _11927_ (
    .A(_03736_),
    .B(_03737_),
    .Y(_03738_)
  );
  OR _11928_ (
    .A(\data_i[5] ),
    .B(_01492_),
    .Y(_03739_)
  );
  AND _11929_ (
    .A(MemWrite_i),
    .B(_03739_),
    .Y(_03740_)
  );
  NAND _11930_ (
    .A(_03738_),
    .B(_03740_),
    .Y(_03741_)
  );
  NAND _11931_ (
    .A(_03728_),
    .B(_03741_),
    .Y(_00189_)
  );
  NAND _11932_ (
    .A(\memory[30][6] ),
    .B(_05361_),
    .Y(_03742_)
  );
  OR _11933_ (
    .A(\memory[30][6] ),
    .B(_01563_),
    .Y(_03743_)
  );
  OR _11934_ (
    .A(\data_i[30] ),
    .B(_01564_),
    .Y(_03744_)
  );
  NAND _11935_ (
    .A(_03743_),
    .B(_03744_),
    .Y(_03745_)
  );
  NAND _11936_ (
    .A(_01463_),
    .B(_03745_),
    .Y(_03746_)
  );
  OR _11937_ (
    .A(\data_i[22] ),
    .B(_01463_),
    .Y(_03747_)
  );
  AND _11938_ (
    .A(_03746_),
    .B(_03747_),
    .Y(_03748_)
  );
  NAND _11939_ (
    .A(\data_i[14] ),
    .B(_01510_),
    .Y(_03749_)
  );
  AND _11940_ (
    .A(_01492_),
    .B(_03749_),
    .Y(_03750_)
  );
  NAND _11941_ (
    .A(_01511_),
    .B(_03748_),
    .Y(_03751_)
  );
  NAND _11942_ (
    .A(_03750_),
    .B(_03751_),
    .Y(_03752_)
  );
  OR _11943_ (
    .A(\data_i[6] ),
    .B(_01492_),
    .Y(_03753_)
  );
  AND _11944_ (
    .A(MemWrite_i),
    .B(_03753_),
    .Y(_03754_)
  );
  NAND _11945_ (
    .A(_03752_),
    .B(_03754_),
    .Y(_03755_)
  );
  NAND _11946_ (
    .A(_03742_),
    .B(_03755_),
    .Y(_00190_)
  );
  NAND _11947_ (
    .A(\memory[30][7] ),
    .B(_05361_),
    .Y(_03756_)
  );
  OR _11948_ (
    .A(\memory[30][7] ),
    .B(_01563_),
    .Y(_03757_)
  );
  OR _11949_ (
    .A(\data_i[31] ),
    .B(_01564_),
    .Y(_03758_)
  );
  NAND _11950_ (
    .A(_03757_),
    .B(_03758_),
    .Y(_03759_)
  );
  NAND _11951_ (
    .A(_01463_),
    .B(_03759_),
    .Y(_03760_)
  );
  OR _11952_ (
    .A(\data_i[23] ),
    .B(_01463_),
    .Y(_03761_)
  );
  AND _11953_ (
    .A(_03760_),
    .B(_03761_),
    .Y(_03762_)
  );
  NAND _11954_ (
    .A(\data_i[15] ),
    .B(_01510_),
    .Y(_03763_)
  );
  AND _11955_ (
    .A(_01492_),
    .B(_03763_),
    .Y(_03764_)
  );
  NAND _11956_ (
    .A(_01511_),
    .B(_03762_),
    .Y(_03765_)
  );
  NAND _11957_ (
    .A(_03764_),
    .B(_03765_),
    .Y(_03766_)
  );
  OR _11958_ (
    .A(\data_i[7] ),
    .B(_01492_),
    .Y(_03767_)
  );
  AND _11959_ (
    .A(MemWrite_i),
    .B(_03767_),
    .Y(_03768_)
  );
  NAND _11960_ (
    .A(_03766_),
    .B(_03768_),
    .Y(_03769_)
  );
  NAND _11961_ (
    .A(_03756_),
    .B(_03769_),
    .Y(_00191_)
  );
  NAND _11962_ (
    .A(\memory[29][0] ),
    .B(_05361_),
    .Y(_03770_)
  );
  OR _11963_ (
    .A(\memory[29][0] ),
    .B(_01484_),
    .Y(_03771_)
  );
  OR _11964_ (
    .A(\data_i[24] ),
    .B(_01485_),
    .Y(_03772_)
  );
  NAND _11965_ (
    .A(_03771_),
    .B(_03772_),
    .Y(_03773_)
  );
  NAND _11966_ (
    .A(_01564_),
    .B(_03773_),
    .Y(_03774_)
  );
  OR _11967_ (
    .A(\data_i[16] ),
    .B(_01564_),
    .Y(_03775_)
  );
  AND _11968_ (
    .A(_03774_),
    .B(_03775_),
    .Y(_03776_)
  );
  NAND _11969_ (
    .A(\data_i[8] ),
    .B(_01462_),
    .Y(_03777_)
  );
  AND _11970_ (
    .A(_01511_),
    .B(_03777_),
    .Y(_03778_)
  );
  NAND _11971_ (
    .A(_01463_),
    .B(_03776_),
    .Y(_03779_)
  );
  NAND _11972_ (
    .A(_03778_),
    .B(_03779_),
    .Y(_03780_)
  );
  OR _11973_ (
    .A(\data_i[0] ),
    .B(_01511_),
    .Y(_03781_)
  );
  AND _11974_ (
    .A(MemWrite_i),
    .B(_03781_),
    .Y(_03782_)
  );
  NAND _11975_ (
    .A(_03780_),
    .B(_03782_),
    .Y(_03783_)
  );
  NAND _11976_ (
    .A(_03770_),
    .B(_03783_),
    .Y(_00168_)
  );
  OR _11977_ (
    .A(\memory[29][1] ),
    .B(MemWrite_i),
    .Y(_03784_)
  );
  NAND _11978_ (
    .A(\data_i[25] ),
    .B(_01484_),
    .Y(_03785_)
  );
  NAND _11979_ (
    .A(\memory[29][1] ),
    .B(_01485_),
    .Y(_03786_)
  );
  NAND _11980_ (
    .A(_03785_),
    .B(_03786_),
    .Y(_03787_)
  );
  NAND _11981_ (
    .A(_01564_),
    .B(_03787_),
    .Y(_03788_)
  );
  NAND _11982_ (
    .A(\data_i[17] ),
    .B(_01563_),
    .Y(_03789_)
  );
  AND _11983_ (
    .A(_01463_),
    .B(_03789_),
    .Y(_03790_)
  );
  NAND _11984_ (
    .A(_03788_),
    .B(_03790_),
    .Y(_03791_)
  );
  OR _11985_ (
    .A(\data_i[9] ),
    .B(_01463_),
    .Y(_03792_)
  );
  AND _11986_ (
    .A(_01511_),
    .B(_03792_),
    .Y(_03793_)
  );
  NAND _11987_ (
    .A(_03791_),
    .B(_03793_),
    .Y(_03794_)
  );
  NAND _11988_ (
    .A(\data_i[1] ),
    .B(_01510_),
    .Y(_03795_)
  );
  AND _11989_ (
    .A(MemWrite_i),
    .B(_03795_),
    .Y(_03796_)
  );
  NAND _11990_ (
    .A(_03794_),
    .B(_03796_),
    .Y(_03797_)
  );
  AND _11991_ (
    .A(_03784_),
    .B(_03797_),
    .Y(_00169_)
  );
  NAND _11992_ (
    .A(\memory[29][2] ),
    .B(_05361_),
    .Y(_03798_)
  );
  OR _11993_ (
    .A(\memory[29][2] ),
    .B(_01484_),
    .Y(_03799_)
  );
  OR _11994_ (
    .A(\data_i[26] ),
    .B(_01485_),
    .Y(_03800_)
  );
  NAND _11995_ (
    .A(_03799_),
    .B(_03800_),
    .Y(_03801_)
  );
  NAND _11996_ (
    .A(_01564_),
    .B(_03801_),
    .Y(_03802_)
  );
  OR _11997_ (
    .A(\data_i[18] ),
    .B(_01564_),
    .Y(_03803_)
  );
  AND _11998_ (
    .A(_03802_),
    .B(_03803_),
    .Y(_03804_)
  );
  NAND _11999_ (
    .A(\data_i[10] ),
    .B(_01462_),
    .Y(_03805_)
  );
  AND _12000_ (
    .A(_01511_),
    .B(_03805_),
    .Y(_03806_)
  );
  NAND _12001_ (
    .A(_01463_),
    .B(_03804_),
    .Y(_03807_)
  );
  NAND _12002_ (
    .A(_03806_),
    .B(_03807_),
    .Y(_03808_)
  );
  OR _12003_ (
    .A(\data_i[2] ),
    .B(_01511_),
    .Y(_03809_)
  );
  AND _12004_ (
    .A(MemWrite_i),
    .B(_03809_),
    .Y(_03810_)
  );
  NAND _12005_ (
    .A(_03808_),
    .B(_03810_),
    .Y(_03811_)
  );
  NAND _12006_ (
    .A(_03798_),
    .B(_03811_),
    .Y(_00170_)
  );
  NAND _12007_ (
    .A(\memory[29][3] ),
    .B(_05361_),
    .Y(_03812_)
  );
  OR _12008_ (
    .A(\memory[29][3] ),
    .B(_01484_),
    .Y(_03813_)
  );
  OR _12009_ (
    .A(\data_i[27] ),
    .B(_01485_),
    .Y(_03814_)
  );
  NAND _12010_ (
    .A(_03813_),
    .B(_03814_),
    .Y(_03815_)
  );
  NAND _12011_ (
    .A(_01564_),
    .B(_03815_),
    .Y(_03816_)
  );
  OR _12012_ (
    .A(\data_i[19] ),
    .B(_01564_),
    .Y(_03817_)
  );
  AND _12013_ (
    .A(_03816_),
    .B(_03817_),
    .Y(_03818_)
  );
  NAND _12014_ (
    .A(\data_i[11] ),
    .B(_01462_),
    .Y(_03819_)
  );
  AND _12015_ (
    .A(_01511_),
    .B(_03819_),
    .Y(_03820_)
  );
  NAND _12016_ (
    .A(_01463_),
    .B(_03818_),
    .Y(_03821_)
  );
  NAND _12017_ (
    .A(_03820_),
    .B(_03821_),
    .Y(_03822_)
  );
  OR _12018_ (
    .A(\data_i[3] ),
    .B(_01511_),
    .Y(_03823_)
  );
  AND _12019_ (
    .A(MemWrite_i),
    .B(_03823_),
    .Y(_03824_)
  );
  NAND _12020_ (
    .A(_03822_),
    .B(_03824_),
    .Y(_03825_)
  );
  NAND _12021_ (
    .A(_03812_),
    .B(_03825_),
    .Y(_00171_)
  );
  NAND _12022_ (
    .A(\memory[29][4] ),
    .B(_05361_),
    .Y(_03826_)
  );
  OR _12023_ (
    .A(\memory[29][4] ),
    .B(_01484_),
    .Y(_03827_)
  );
  OR _12024_ (
    .A(\data_i[28] ),
    .B(_01485_),
    .Y(_03828_)
  );
  NAND _12025_ (
    .A(_03827_),
    .B(_03828_),
    .Y(_03829_)
  );
  NAND _12026_ (
    .A(_01564_),
    .B(_03829_),
    .Y(_03830_)
  );
  OR _12027_ (
    .A(\data_i[20] ),
    .B(_01564_),
    .Y(_03831_)
  );
  AND _12028_ (
    .A(_03830_),
    .B(_03831_),
    .Y(_03832_)
  );
  NAND _12029_ (
    .A(\data_i[12] ),
    .B(_01462_),
    .Y(_03833_)
  );
  AND _12030_ (
    .A(_01511_),
    .B(_03833_),
    .Y(_03834_)
  );
  NAND _12031_ (
    .A(_01463_),
    .B(_03832_),
    .Y(_03835_)
  );
  NAND _12032_ (
    .A(_03834_),
    .B(_03835_),
    .Y(_03836_)
  );
  OR _12033_ (
    .A(\data_i[4] ),
    .B(_01511_),
    .Y(_03837_)
  );
  AND _12034_ (
    .A(MemWrite_i),
    .B(_03837_),
    .Y(_03838_)
  );
  NAND _12035_ (
    .A(_03836_),
    .B(_03838_),
    .Y(_03839_)
  );
  NAND _12036_ (
    .A(_03826_),
    .B(_03839_),
    .Y(_00172_)
  );
  NAND _12037_ (
    .A(\memory[29][5] ),
    .B(_05361_),
    .Y(_03840_)
  );
  OR _12038_ (
    .A(\memory[29][5] ),
    .B(_01484_),
    .Y(_03841_)
  );
  OR _12039_ (
    .A(\data_i[29] ),
    .B(_01485_),
    .Y(_03842_)
  );
  NAND _12040_ (
    .A(_03841_),
    .B(_03842_),
    .Y(_03843_)
  );
  NAND _12041_ (
    .A(_01564_),
    .B(_03843_),
    .Y(_03844_)
  );
  OR _12042_ (
    .A(\data_i[21] ),
    .B(_01564_),
    .Y(_03845_)
  );
  AND _12043_ (
    .A(_03844_),
    .B(_03845_),
    .Y(_03846_)
  );
  NAND _12044_ (
    .A(\data_i[13] ),
    .B(_01462_),
    .Y(_03847_)
  );
  AND _12045_ (
    .A(_01511_),
    .B(_03847_),
    .Y(_03848_)
  );
  NAND _12046_ (
    .A(_01463_),
    .B(_03846_),
    .Y(_03849_)
  );
  NAND _12047_ (
    .A(_03848_),
    .B(_03849_),
    .Y(_03850_)
  );
  OR _12048_ (
    .A(\data_i[5] ),
    .B(_01511_),
    .Y(_03851_)
  );
  AND _12049_ (
    .A(MemWrite_i),
    .B(_03851_),
    .Y(_03852_)
  );
  NAND _12050_ (
    .A(_03850_),
    .B(_03852_),
    .Y(_03853_)
  );
  NAND _12051_ (
    .A(_03840_),
    .B(_03853_),
    .Y(_00173_)
  );
  NAND _12052_ (
    .A(\memory[29][6] ),
    .B(_05361_),
    .Y(_03854_)
  );
  OR _12053_ (
    .A(\memory[29][6] ),
    .B(_01484_),
    .Y(_03855_)
  );
  OR _12054_ (
    .A(\data_i[30] ),
    .B(_01485_),
    .Y(_03856_)
  );
  NAND _12055_ (
    .A(_03855_),
    .B(_03856_),
    .Y(_03857_)
  );
  NAND _12056_ (
    .A(_01564_),
    .B(_03857_),
    .Y(_03858_)
  );
  OR _12057_ (
    .A(\data_i[22] ),
    .B(_01564_),
    .Y(_03859_)
  );
  AND _12058_ (
    .A(_03858_),
    .B(_03859_),
    .Y(_03860_)
  );
  NAND _12059_ (
    .A(\data_i[14] ),
    .B(_01462_),
    .Y(_03861_)
  );
  AND _12060_ (
    .A(_01511_),
    .B(_03861_),
    .Y(_03862_)
  );
  NAND _12061_ (
    .A(_01463_),
    .B(_03860_),
    .Y(_03863_)
  );
  NAND _12062_ (
    .A(_03862_),
    .B(_03863_),
    .Y(_03864_)
  );
  OR _12063_ (
    .A(\data_i[6] ),
    .B(_01511_),
    .Y(_03865_)
  );
  AND _12064_ (
    .A(MemWrite_i),
    .B(_03865_),
    .Y(_03866_)
  );
  NAND _12065_ (
    .A(_03864_),
    .B(_03866_),
    .Y(_03867_)
  );
  NAND _12066_ (
    .A(_03854_),
    .B(_03867_),
    .Y(_00174_)
  );
  NAND _12067_ (
    .A(\memory[29][7] ),
    .B(_05361_),
    .Y(_03868_)
  );
  OR _12068_ (
    .A(\memory[29][7] ),
    .B(_01484_),
    .Y(_03869_)
  );
  OR _12069_ (
    .A(\data_i[31] ),
    .B(_01485_),
    .Y(_03870_)
  );
  NAND _12070_ (
    .A(_03869_),
    .B(_03870_),
    .Y(_03871_)
  );
  NAND _12071_ (
    .A(_01564_),
    .B(_03871_),
    .Y(_03872_)
  );
  OR _12072_ (
    .A(\data_i[23] ),
    .B(_01564_),
    .Y(_03873_)
  );
  AND _12073_ (
    .A(_03872_),
    .B(_03873_),
    .Y(_03874_)
  );
  NAND _12074_ (
    .A(\data_i[15] ),
    .B(_01462_),
    .Y(_03875_)
  );
  AND _12075_ (
    .A(_01511_),
    .B(_03875_),
    .Y(_03876_)
  );
  NAND _12076_ (
    .A(_01463_),
    .B(_03874_),
    .Y(_03877_)
  );
  NAND _12077_ (
    .A(_03876_),
    .B(_03877_),
    .Y(_03878_)
  );
  OR _12078_ (
    .A(\data_i[7] ),
    .B(_01511_),
    .Y(_03879_)
  );
  AND _12079_ (
    .A(MemWrite_i),
    .B(_03879_),
    .Y(_03880_)
  );
  NAND _12080_ (
    .A(_03878_),
    .B(_03880_),
    .Y(_03881_)
  );
  NAND _12081_ (
    .A(_03868_),
    .B(_03881_),
    .Y(_00175_)
  );
  NAND _12082_ (
    .A(\memory[28][0] ),
    .B(_05361_),
    .Y(_03882_)
  );
  OR _12083_ (
    .A(\memory[28][0] ),
    .B(_01559_),
    .Y(_03883_)
  );
  OR _12084_ (
    .A(\data_i[24] ),
    .B(_01560_),
    .Y(_03884_)
  );
  NAND _12085_ (
    .A(_03883_),
    .B(_03884_),
    .Y(_03885_)
  );
  NAND _12086_ (
    .A(_01485_),
    .B(_03885_),
    .Y(_03886_)
  );
  OR _12087_ (
    .A(\data_i[16] ),
    .B(_01485_),
    .Y(_03887_)
  );
  AND _12088_ (
    .A(_03886_),
    .B(_03887_),
    .Y(_03888_)
  );
  NAND _12089_ (
    .A(\data_i[8] ),
    .B(_01563_),
    .Y(_03889_)
  );
  AND _12090_ (
    .A(_01463_),
    .B(_03889_),
    .Y(_03890_)
  );
  NAND _12091_ (
    .A(_01564_),
    .B(_03888_),
    .Y(_03891_)
  );
  NAND _12092_ (
    .A(_03890_),
    .B(_03891_),
    .Y(_03892_)
  );
  OR _12093_ (
    .A(\data_i[0] ),
    .B(_01463_),
    .Y(_03893_)
  );
  AND _12094_ (
    .A(MemWrite_i),
    .B(_03893_),
    .Y(_03894_)
  );
  NAND _12095_ (
    .A(_03892_),
    .B(_03894_),
    .Y(_03895_)
  );
  NAND _12096_ (
    .A(_03882_),
    .B(_03895_),
    .Y(_00160_)
  );
  NAND _12097_ (
    .A(\memory[28][1] ),
    .B(_05361_),
    .Y(_03896_)
  );
  OR _12098_ (
    .A(\memory[28][1] ),
    .B(_01559_),
    .Y(_03897_)
  );
  OR _12099_ (
    .A(\data_i[25] ),
    .B(_01560_),
    .Y(_03898_)
  );
  NAND _12100_ (
    .A(_03897_),
    .B(_03898_),
    .Y(_03899_)
  );
  NAND _12101_ (
    .A(_01485_),
    .B(_03899_),
    .Y(_03900_)
  );
  OR _12102_ (
    .A(\data_i[17] ),
    .B(_01485_),
    .Y(_03901_)
  );
  AND _12103_ (
    .A(_03900_),
    .B(_03901_),
    .Y(_03902_)
  );
  NAND _12104_ (
    .A(\data_i[9] ),
    .B(_01563_),
    .Y(_03903_)
  );
  AND _12105_ (
    .A(_01463_),
    .B(_03903_),
    .Y(_03904_)
  );
  NAND _12106_ (
    .A(_01564_),
    .B(_03902_),
    .Y(_03905_)
  );
  NAND _12107_ (
    .A(_03904_),
    .B(_03905_),
    .Y(_03906_)
  );
  OR _12108_ (
    .A(\data_i[1] ),
    .B(_01463_),
    .Y(_03907_)
  );
  AND _12109_ (
    .A(MemWrite_i),
    .B(_03907_),
    .Y(_03908_)
  );
  NAND _12110_ (
    .A(_03906_),
    .B(_03908_),
    .Y(_03909_)
  );
  NAND _12111_ (
    .A(_03896_),
    .B(_03909_),
    .Y(_00161_)
  );
  NAND _12112_ (
    .A(\memory[28][2] ),
    .B(_05361_),
    .Y(_03910_)
  );
  OR _12113_ (
    .A(\memory[28][2] ),
    .B(_01559_),
    .Y(_03911_)
  );
  OR _12114_ (
    .A(\data_i[26] ),
    .B(_01560_),
    .Y(_03912_)
  );
  NAND _12115_ (
    .A(_03911_),
    .B(_03912_),
    .Y(_03913_)
  );
  NAND _12116_ (
    .A(_01485_),
    .B(_03913_),
    .Y(_03914_)
  );
  OR _12117_ (
    .A(\data_i[18] ),
    .B(_01485_),
    .Y(_03915_)
  );
  AND _12118_ (
    .A(_03914_),
    .B(_03915_),
    .Y(_03916_)
  );
  NAND _12119_ (
    .A(\data_i[10] ),
    .B(_01563_),
    .Y(_03917_)
  );
  AND _12120_ (
    .A(_01463_),
    .B(_03917_),
    .Y(_03918_)
  );
  NAND _12121_ (
    .A(_01564_),
    .B(_03916_),
    .Y(_03919_)
  );
  NAND _12122_ (
    .A(_03918_),
    .B(_03919_),
    .Y(_03920_)
  );
  OR _12123_ (
    .A(\data_i[2] ),
    .B(_01463_),
    .Y(_03921_)
  );
  AND _12124_ (
    .A(MemWrite_i),
    .B(_03921_),
    .Y(_03922_)
  );
  NAND _12125_ (
    .A(_03920_),
    .B(_03922_),
    .Y(_03923_)
  );
  NAND _12126_ (
    .A(_03910_),
    .B(_03923_),
    .Y(_00162_)
  );
  NAND _12127_ (
    .A(\memory[28][3] ),
    .B(_05361_),
    .Y(_03924_)
  );
  OR _12128_ (
    .A(\memory[28][3] ),
    .B(_01559_),
    .Y(_03925_)
  );
  OR _12129_ (
    .A(\data_i[27] ),
    .B(_01560_),
    .Y(_03926_)
  );
  NAND _12130_ (
    .A(_03925_),
    .B(_03926_),
    .Y(_03927_)
  );
  NAND _12131_ (
    .A(_01485_),
    .B(_03927_),
    .Y(_03928_)
  );
  OR _12132_ (
    .A(\data_i[19] ),
    .B(_01485_),
    .Y(_03929_)
  );
  AND _12133_ (
    .A(_03928_),
    .B(_03929_),
    .Y(_03930_)
  );
  NAND _12134_ (
    .A(\data_i[11] ),
    .B(_01563_),
    .Y(_03931_)
  );
  AND _12135_ (
    .A(_01463_),
    .B(_03931_),
    .Y(_03932_)
  );
  NAND _12136_ (
    .A(_01564_),
    .B(_03930_),
    .Y(_03933_)
  );
  NAND _12137_ (
    .A(_03932_),
    .B(_03933_),
    .Y(_03934_)
  );
  OR _12138_ (
    .A(\data_i[3] ),
    .B(_01463_),
    .Y(_03935_)
  );
  AND _12139_ (
    .A(MemWrite_i),
    .B(_03935_),
    .Y(_03936_)
  );
  NAND _12140_ (
    .A(_03934_),
    .B(_03936_),
    .Y(_03937_)
  );
  NAND _12141_ (
    .A(_03924_),
    .B(_03937_),
    .Y(_00163_)
  );
  NAND _12142_ (
    .A(\memory[28][4] ),
    .B(_05361_),
    .Y(_03938_)
  );
  OR _12143_ (
    .A(\memory[28][4] ),
    .B(_01559_),
    .Y(_03939_)
  );
  OR _12144_ (
    .A(\data_i[28] ),
    .B(_01560_),
    .Y(_03940_)
  );
  NAND _12145_ (
    .A(_03939_),
    .B(_03940_),
    .Y(_03941_)
  );
  NAND _12146_ (
    .A(_01485_),
    .B(_03941_),
    .Y(_03942_)
  );
  OR _12147_ (
    .A(\data_i[20] ),
    .B(_01485_),
    .Y(_03943_)
  );
  AND _12148_ (
    .A(_03942_),
    .B(_03943_),
    .Y(_03944_)
  );
  NAND _12149_ (
    .A(\data_i[12] ),
    .B(_01563_),
    .Y(_03945_)
  );
  AND _12150_ (
    .A(_01463_),
    .B(_03945_),
    .Y(_03946_)
  );
  NAND _12151_ (
    .A(_01564_),
    .B(_03944_),
    .Y(_03947_)
  );
  NAND _12152_ (
    .A(_03946_),
    .B(_03947_),
    .Y(_03948_)
  );
  OR _12153_ (
    .A(\data_i[4] ),
    .B(_01463_),
    .Y(_03949_)
  );
  AND _12154_ (
    .A(MemWrite_i),
    .B(_03949_),
    .Y(_03950_)
  );
  NAND _12155_ (
    .A(_03948_),
    .B(_03950_),
    .Y(_03951_)
  );
  NAND _12156_ (
    .A(_03938_),
    .B(_03951_),
    .Y(_00164_)
  );
  NAND _12157_ (
    .A(\memory[28][5] ),
    .B(_05361_),
    .Y(_03952_)
  );
  OR _12158_ (
    .A(\memory[28][5] ),
    .B(_01559_),
    .Y(_03953_)
  );
  OR _12159_ (
    .A(\data_i[29] ),
    .B(_01560_),
    .Y(_03954_)
  );
  NAND _12160_ (
    .A(_03953_),
    .B(_03954_),
    .Y(_03955_)
  );
  NAND _12161_ (
    .A(_01485_),
    .B(_03955_),
    .Y(_03956_)
  );
  OR _12162_ (
    .A(\data_i[21] ),
    .B(_01485_),
    .Y(_03957_)
  );
  AND _12163_ (
    .A(_03956_),
    .B(_03957_),
    .Y(_03958_)
  );
  NAND _12164_ (
    .A(_01564_),
    .B(_03958_),
    .Y(_03959_)
  );
  NAND _12165_ (
    .A(\data_i[13] ),
    .B(_01563_),
    .Y(_03960_)
  );
  AND _12166_ (
    .A(_01463_),
    .B(_03960_),
    .Y(_03961_)
  );
  NAND _12167_ (
    .A(_03959_),
    .B(_03961_),
    .Y(_03962_)
  );
  OR _12168_ (
    .A(\data_i[5] ),
    .B(_01463_),
    .Y(_03963_)
  );
  AND _12169_ (
    .A(MemWrite_i),
    .B(_03963_),
    .Y(_03964_)
  );
  NAND _12170_ (
    .A(_03962_),
    .B(_03964_),
    .Y(_03965_)
  );
  NAND _12171_ (
    .A(_03952_),
    .B(_03965_),
    .Y(_00165_)
  );
  NAND _12172_ (
    .A(\memory[28][6] ),
    .B(_05361_),
    .Y(_03966_)
  );
  OR _12173_ (
    .A(\memory[28][6] ),
    .B(_01559_),
    .Y(_03967_)
  );
  OR _12174_ (
    .A(\data_i[30] ),
    .B(_01560_),
    .Y(_03968_)
  );
  NAND _12175_ (
    .A(_03967_),
    .B(_03968_),
    .Y(_03969_)
  );
  NAND _12176_ (
    .A(_01485_),
    .B(_03969_),
    .Y(_03970_)
  );
  OR _12177_ (
    .A(\data_i[22] ),
    .B(_01485_),
    .Y(_03971_)
  );
  AND _12178_ (
    .A(_03970_),
    .B(_03971_),
    .Y(_03972_)
  );
  NAND _12179_ (
    .A(\data_i[14] ),
    .B(_01563_),
    .Y(_03973_)
  );
  AND _12180_ (
    .A(_01463_),
    .B(_03973_),
    .Y(_03974_)
  );
  NAND _12181_ (
    .A(_01564_),
    .B(_03972_),
    .Y(_03975_)
  );
  NAND _12182_ (
    .A(_03974_),
    .B(_03975_),
    .Y(_03976_)
  );
  OR _12183_ (
    .A(\data_i[6] ),
    .B(_01463_),
    .Y(_03977_)
  );
  AND _12184_ (
    .A(MemWrite_i),
    .B(_03977_),
    .Y(_03978_)
  );
  NAND _12185_ (
    .A(_03976_),
    .B(_03978_),
    .Y(_03979_)
  );
  NAND _12186_ (
    .A(_03966_),
    .B(_03979_),
    .Y(_00166_)
  );
  NAND _12187_ (
    .A(\memory[28][7] ),
    .B(_05361_),
    .Y(_03980_)
  );
  OR _12188_ (
    .A(\memory[28][7] ),
    .B(_01559_),
    .Y(_03981_)
  );
  OR _12189_ (
    .A(\data_i[31] ),
    .B(_01560_),
    .Y(_03982_)
  );
  NAND _12190_ (
    .A(_03981_),
    .B(_03982_),
    .Y(_03983_)
  );
  NAND _12191_ (
    .A(_01485_),
    .B(_03983_),
    .Y(_03984_)
  );
  OR _12192_ (
    .A(\data_i[23] ),
    .B(_01485_),
    .Y(_03985_)
  );
  AND _12193_ (
    .A(_03984_),
    .B(_03985_),
    .Y(_03986_)
  );
  NAND _12194_ (
    .A(\data_i[15] ),
    .B(_01563_),
    .Y(_03987_)
  );
  AND _12195_ (
    .A(_01463_),
    .B(_03987_),
    .Y(_03988_)
  );
  NAND _12196_ (
    .A(_01564_),
    .B(_03986_),
    .Y(_03989_)
  );
  NAND _12197_ (
    .A(_03988_),
    .B(_03989_),
    .Y(_03990_)
  );
  OR _12198_ (
    .A(\data_i[7] ),
    .B(_01463_),
    .Y(_03991_)
  );
  AND _12199_ (
    .A(MemWrite_i),
    .B(_03991_),
    .Y(_03992_)
  );
  NAND _12200_ (
    .A(_03990_),
    .B(_03992_),
    .Y(_03993_)
  );
  NAND _12201_ (
    .A(_03980_),
    .B(_03993_),
    .Y(_00167_)
  );
  OR _12202_ (
    .A(\memory[27][0] ),
    .B(MemWrite_i),
    .Y(_03994_)
  );
  NAND _12203_ (
    .A(\data_i[24] ),
    .B(_01550_),
    .Y(_03995_)
  );
  NAND _12204_ (
    .A(\memory[27][0] ),
    .B(_01551_),
    .Y(_03996_)
  );
  NAND _12205_ (
    .A(_03995_),
    .B(_03996_),
    .Y(_03997_)
  );
  NAND _12206_ (
    .A(_01560_),
    .B(_03997_),
    .Y(_03998_)
  );
  NAND _12207_ (
    .A(\data_i[16] ),
    .B(_01559_),
    .Y(_03999_)
  );
  AND _12208_ (
    .A(_01485_),
    .B(_03999_),
    .Y(_04000_)
  );
  NAND _12209_ (
    .A(_03998_),
    .B(_04000_),
    .Y(_04001_)
  );
  OR _12210_ (
    .A(\data_i[8] ),
    .B(_01485_),
    .Y(_04002_)
  );
  AND _12211_ (
    .A(_01564_),
    .B(_04002_),
    .Y(_04003_)
  );
  NAND _12212_ (
    .A(_04001_),
    .B(_04003_),
    .Y(_04004_)
  );
  NAND _12213_ (
    .A(\data_i[0] ),
    .B(_01563_),
    .Y(_04005_)
  );
  AND _12214_ (
    .A(MemWrite_i),
    .B(_04005_),
    .Y(_04006_)
  );
  NAND _12215_ (
    .A(_04004_),
    .B(_04006_),
    .Y(_04007_)
  );
  AND _12216_ (
    .A(_03994_),
    .B(_04007_),
    .Y(_00152_)
  );
  NAND _12217_ (
    .A(\memory[27][1] ),
    .B(_05361_),
    .Y(_04008_)
  );
  OR _12218_ (
    .A(\memory[27][1] ),
    .B(_01550_),
    .Y(_04009_)
  );
  OR _12219_ (
    .A(\data_i[25] ),
    .B(_01551_),
    .Y(_04010_)
  );
  NAND _12220_ (
    .A(_04009_),
    .B(_04010_),
    .Y(_04011_)
  );
  NAND _12221_ (
    .A(_01560_),
    .B(_04011_),
    .Y(_04012_)
  );
  OR _12222_ (
    .A(\data_i[17] ),
    .B(_01560_),
    .Y(_04013_)
  );
  AND _12223_ (
    .A(_04012_),
    .B(_04013_),
    .Y(_04014_)
  );
  NAND _12224_ (
    .A(\data_i[9] ),
    .B(_01484_),
    .Y(_04015_)
  );
  AND _12225_ (
    .A(_01564_),
    .B(_04015_),
    .Y(_04016_)
  );
  NAND _12226_ (
    .A(_01485_),
    .B(_04014_),
    .Y(_04017_)
  );
  NAND _12227_ (
    .A(_04016_),
    .B(_04017_),
    .Y(_04018_)
  );
  OR _12228_ (
    .A(\data_i[1] ),
    .B(_01564_),
    .Y(_04019_)
  );
  AND _12229_ (
    .A(MemWrite_i),
    .B(_04019_),
    .Y(_04020_)
  );
  NAND _12230_ (
    .A(_04018_),
    .B(_04020_),
    .Y(_04021_)
  );
  NAND _12231_ (
    .A(_04008_),
    .B(_04021_),
    .Y(_00153_)
  );
  NAND _12232_ (
    .A(\memory[27][2] ),
    .B(_05361_),
    .Y(_04022_)
  );
  OR _12233_ (
    .A(\memory[27][2] ),
    .B(_01550_),
    .Y(_04023_)
  );
  OR _12234_ (
    .A(\data_i[26] ),
    .B(_01551_),
    .Y(_04024_)
  );
  NAND _12235_ (
    .A(_04023_),
    .B(_04024_),
    .Y(_04025_)
  );
  NAND _12236_ (
    .A(_01560_),
    .B(_04025_),
    .Y(_04026_)
  );
  OR _12237_ (
    .A(\data_i[18] ),
    .B(_01560_),
    .Y(_04027_)
  );
  AND _12238_ (
    .A(_04026_),
    .B(_04027_),
    .Y(_04028_)
  );
  NAND _12239_ (
    .A(\data_i[10] ),
    .B(_01484_),
    .Y(_04029_)
  );
  AND _12240_ (
    .A(_01564_),
    .B(_04029_),
    .Y(_04030_)
  );
  NAND _12241_ (
    .A(_01485_),
    .B(_04028_),
    .Y(_04031_)
  );
  NAND _12242_ (
    .A(_04030_),
    .B(_04031_),
    .Y(_04032_)
  );
  OR _12243_ (
    .A(\data_i[2] ),
    .B(_01564_),
    .Y(_04033_)
  );
  AND _12244_ (
    .A(MemWrite_i),
    .B(_04033_),
    .Y(_04034_)
  );
  NAND _12245_ (
    .A(_04032_),
    .B(_04034_),
    .Y(_04035_)
  );
  NAND _12246_ (
    .A(_04022_),
    .B(_04035_),
    .Y(_00154_)
  );
  NAND _12247_ (
    .A(\memory[27][3] ),
    .B(_05361_),
    .Y(_04036_)
  );
  OR _12248_ (
    .A(\memory[27][3] ),
    .B(_01550_),
    .Y(_04037_)
  );
  OR _12249_ (
    .A(\data_i[27] ),
    .B(_01551_),
    .Y(_04038_)
  );
  NAND _12250_ (
    .A(_04037_),
    .B(_04038_),
    .Y(_04039_)
  );
  NAND _12251_ (
    .A(_01560_),
    .B(_04039_),
    .Y(_04040_)
  );
  OR _12252_ (
    .A(\data_i[19] ),
    .B(_01560_),
    .Y(_04041_)
  );
  AND _12253_ (
    .A(_04040_),
    .B(_04041_),
    .Y(_04042_)
  );
  NAND _12254_ (
    .A(\data_i[11] ),
    .B(_01484_),
    .Y(_04043_)
  );
  AND _12255_ (
    .A(_01564_),
    .B(_04043_),
    .Y(_04044_)
  );
  NAND _12256_ (
    .A(_01485_),
    .B(_04042_),
    .Y(_04045_)
  );
  NAND _12257_ (
    .A(_04044_),
    .B(_04045_),
    .Y(_04046_)
  );
  OR _12258_ (
    .A(\data_i[3] ),
    .B(_01564_),
    .Y(_04047_)
  );
  AND _12259_ (
    .A(MemWrite_i),
    .B(_04047_),
    .Y(_04048_)
  );
  NAND _12260_ (
    .A(_04046_),
    .B(_04048_),
    .Y(_04049_)
  );
  NAND _12261_ (
    .A(_04036_),
    .B(_04049_),
    .Y(_00155_)
  );
  NAND _12262_ (
    .A(\memory[27][4] ),
    .B(_05361_),
    .Y(_04050_)
  );
  OR _12263_ (
    .A(\memory[27][4] ),
    .B(_01550_),
    .Y(_04051_)
  );
  OR _12264_ (
    .A(\data_i[28] ),
    .B(_01551_),
    .Y(_04052_)
  );
  NAND _12265_ (
    .A(_04051_),
    .B(_04052_),
    .Y(_04053_)
  );
  NAND _12266_ (
    .A(_01560_),
    .B(_04053_),
    .Y(_04054_)
  );
  OR _12267_ (
    .A(\data_i[20] ),
    .B(_01560_),
    .Y(_04055_)
  );
  AND _12268_ (
    .A(_04054_),
    .B(_04055_),
    .Y(_04056_)
  );
  NAND _12269_ (
    .A(\data_i[12] ),
    .B(_01484_),
    .Y(_04057_)
  );
  AND _12270_ (
    .A(_01564_),
    .B(_04057_),
    .Y(_04058_)
  );
  NAND _12271_ (
    .A(_01485_),
    .B(_04056_),
    .Y(_04059_)
  );
  NAND _12272_ (
    .A(_04058_),
    .B(_04059_),
    .Y(_04060_)
  );
  OR _12273_ (
    .A(\data_i[4] ),
    .B(_01564_),
    .Y(_04061_)
  );
  AND _12274_ (
    .A(MemWrite_i),
    .B(_04061_),
    .Y(_04062_)
  );
  NAND _12275_ (
    .A(_04060_),
    .B(_04062_),
    .Y(_04063_)
  );
  NAND _12276_ (
    .A(_04050_),
    .B(_04063_),
    .Y(_00156_)
  );
  NAND _12277_ (
    .A(\memory[27][5] ),
    .B(_05361_),
    .Y(_04064_)
  );
  OR _12278_ (
    .A(\memory[27][5] ),
    .B(_01550_),
    .Y(_04065_)
  );
  OR _12279_ (
    .A(\data_i[29] ),
    .B(_01551_),
    .Y(_04066_)
  );
  NAND _12280_ (
    .A(_04065_),
    .B(_04066_),
    .Y(_04067_)
  );
  NAND _12281_ (
    .A(_01560_),
    .B(_04067_),
    .Y(_04068_)
  );
  OR _12282_ (
    .A(\data_i[21] ),
    .B(_01560_),
    .Y(_04069_)
  );
  AND _12283_ (
    .A(_04068_),
    .B(_04069_),
    .Y(_04070_)
  );
  NAND _12284_ (
    .A(\data_i[13] ),
    .B(_01484_),
    .Y(_04071_)
  );
  AND _12285_ (
    .A(_01564_),
    .B(_04071_),
    .Y(_04072_)
  );
  NAND _12286_ (
    .A(_01485_),
    .B(_04070_),
    .Y(_04073_)
  );
  NAND _12287_ (
    .A(_04072_),
    .B(_04073_),
    .Y(_04074_)
  );
  OR _12288_ (
    .A(\data_i[5] ),
    .B(_01564_),
    .Y(_04075_)
  );
  AND _12289_ (
    .A(MemWrite_i),
    .B(_04075_),
    .Y(_04076_)
  );
  NAND _12290_ (
    .A(_04074_),
    .B(_04076_),
    .Y(_04077_)
  );
  NAND _12291_ (
    .A(_04064_),
    .B(_04077_),
    .Y(_00157_)
  );
  NAND _12292_ (
    .A(\memory[27][6] ),
    .B(_05361_),
    .Y(_04078_)
  );
  OR _12293_ (
    .A(\memory[27][6] ),
    .B(_01550_),
    .Y(_04079_)
  );
  OR _12294_ (
    .A(\data_i[30] ),
    .B(_01551_),
    .Y(_04080_)
  );
  NAND _12295_ (
    .A(_04079_),
    .B(_04080_),
    .Y(_04081_)
  );
  NAND _12296_ (
    .A(_01560_),
    .B(_04081_),
    .Y(_04082_)
  );
  OR _12297_ (
    .A(\data_i[22] ),
    .B(_01560_),
    .Y(_04083_)
  );
  AND _12298_ (
    .A(_04082_),
    .B(_04083_),
    .Y(_04084_)
  );
  NAND _12299_ (
    .A(\data_i[14] ),
    .B(_01484_),
    .Y(_04085_)
  );
  AND _12300_ (
    .A(_01564_),
    .B(_04085_),
    .Y(_04086_)
  );
  NAND _12301_ (
    .A(_01485_),
    .B(_04084_),
    .Y(_04087_)
  );
  NAND _12302_ (
    .A(_04086_),
    .B(_04087_),
    .Y(_04088_)
  );
  OR _12303_ (
    .A(\data_i[6] ),
    .B(_01564_),
    .Y(_04089_)
  );
  AND _12304_ (
    .A(MemWrite_i),
    .B(_04089_),
    .Y(_04090_)
  );
  NAND _12305_ (
    .A(_04088_),
    .B(_04090_),
    .Y(_04091_)
  );
  NAND _12306_ (
    .A(_04078_),
    .B(_04091_),
    .Y(_00158_)
  );
  NAND _12307_ (
    .A(\memory[27][7] ),
    .B(_05361_),
    .Y(_04092_)
  );
  OR _12308_ (
    .A(\memory[27][7] ),
    .B(_01550_),
    .Y(_04093_)
  );
  OR _12309_ (
    .A(\data_i[31] ),
    .B(_01551_),
    .Y(_04094_)
  );
  NAND _12310_ (
    .A(_04093_),
    .B(_04094_),
    .Y(_04095_)
  );
  NAND _12311_ (
    .A(_01560_),
    .B(_04095_),
    .Y(_04096_)
  );
  OR _12312_ (
    .A(\data_i[23] ),
    .B(_01560_),
    .Y(_04097_)
  );
  AND _12313_ (
    .A(_04096_),
    .B(_04097_),
    .Y(_04098_)
  );
  NAND _12314_ (
    .A(\data_i[15] ),
    .B(_01484_),
    .Y(_04099_)
  );
  AND _12315_ (
    .A(_01564_),
    .B(_04099_),
    .Y(_04100_)
  );
  NAND _12316_ (
    .A(_01485_),
    .B(_04098_),
    .Y(_04101_)
  );
  NAND _12317_ (
    .A(_04100_),
    .B(_04101_),
    .Y(_04102_)
  );
  OR _12318_ (
    .A(\data_i[7] ),
    .B(_01564_),
    .Y(_04103_)
  );
  AND _12319_ (
    .A(MemWrite_i),
    .B(_04103_),
    .Y(_04104_)
  );
  NAND _12320_ (
    .A(_04102_),
    .B(_04104_),
    .Y(_04105_)
  );
  NAND _12321_ (
    .A(_04092_),
    .B(_04105_),
    .Y(_00159_)
  );
  NAND _12322_ (
    .A(\memory[26][0] ),
    .B(_05361_),
    .Y(_04106_)
  );
  OR _12323_ (
    .A(\memory[26][0] ),
    .B(_01546_),
    .Y(_04107_)
  );
  OR _12324_ (
    .A(\data_i[24] ),
    .B(_01547_),
    .Y(_04108_)
  );
  NAND _12325_ (
    .A(_04107_),
    .B(_04108_),
    .Y(_04109_)
  );
  NAND _12326_ (
    .A(_01551_),
    .B(_04109_),
    .Y(_04110_)
  );
  OR _12327_ (
    .A(\data_i[16] ),
    .B(_01551_),
    .Y(_04111_)
  );
  AND _12328_ (
    .A(_04110_),
    .B(_04111_),
    .Y(_04112_)
  );
  NAND _12329_ (
    .A(\data_i[8] ),
    .B(_01559_),
    .Y(_04113_)
  );
  AND _12330_ (
    .A(_01485_),
    .B(_04113_),
    .Y(_04114_)
  );
  NAND _12331_ (
    .A(_01560_),
    .B(_04112_),
    .Y(_04115_)
  );
  NAND _12332_ (
    .A(_04114_),
    .B(_04115_),
    .Y(_04116_)
  );
  OR _12333_ (
    .A(\data_i[0] ),
    .B(_01485_),
    .Y(_04117_)
  );
  AND _12334_ (
    .A(MemWrite_i),
    .B(_04117_),
    .Y(_04118_)
  );
  NAND _12335_ (
    .A(_04116_),
    .B(_04118_),
    .Y(_04119_)
  );
  NAND _12336_ (
    .A(_04106_),
    .B(_04119_),
    .Y(_00144_)
  );
  NAND _12337_ (
    .A(\memory[26][1] ),
    .B(_05361_),
    .Y(_04120_)
  );
  OR _12338_ (
    .A(\memory[26][1] ),
    .B(_01546_),
    .Y(_04121_)
  );
  OR _12339_ (
    .A(\data_i[25] ),
    .B(_01547_),
    .Y(_04122_)
  );
  NAND _12340_ (
    .A(_04121_),
    .B(_04122_),
    .Y(_04123_)
  );
  NAND _12341_ (
    .A(_01551_),
    .B(_04123_),
    .Y(_04124_)
  );
  OR _12342_ (
    .A(\data_i[17] ),
    .B(_01551_),
    .Y(_04125_)
  );
  AND _12343_ (
    .A(_04124_),
    .B(_04125_),
    .Y(_04126_)
  );
  NAND _12344_ (
    .A(\data_i[9] ),
    .B(_01559_),
    .Y(_04127_)
  );
  AND _12345_ (
    .A(_01485_),
    .B(_04127_),
    .Y(_04128_)
  );
  NAND _12346_ (
    .A(_01560_),
    .B(_04126_),
    .Y(_04129_)
  );
  NAND _12347_ (
    .A(_04128_),
    .B(_04129_),
    .Y(_04130_)
  );
  OR _12348_ (
    .A(\data_i[1] ),
    .B(_01485_),
    .Y(_04131_)
  );
  AND _12349_ (
    .A(MemWrite_i),
    .B(_04131_),
    .Y(_04132_)
  );
  NAND _12350_ (
    .A(_04130_),
    .B(_04132_),
    .Y(_04133_)
  );
  NAND _12351_ (
    .A(_04120_),
    .B(_04133_),
    .Y(_00145_)
  );
  NAND _12352_ (
    .A(\memory[26][2] ),
    .B(_05361_),
    .Y(_04134_)
  );
  OR _12353_ (
    .A(\memory[26][2] ),
    .B(_01546_),
    .Y(_04135_)
  );
  OR _12354_ (
    .A(\data_i[26] ),
    .B(_01547_),
    .Y(_04136_)
  );
  NAND _12355_ (
    .A(_04135_),
    .B(_04136_),
    .Y(_04137_)
  );
  NAND _12356_ (
    .A(_01551_),
    .B(_04137_),
    .Y(_04138_)
  );
  OR _12357_ (
    .A(\data_i[18] ),
    .B(_01551_),
    .Y(_04139_)
  );
  AND _12358_ (
    .A(_04138_),
    .B(_04139_),
    .Y(_04140_)
  );
  NAND _12359_ (
    .A(\data_i[10] ),
    .B(_01559_),
    .Y(_04141_)
  );
  AND _12360_ (
    .A(_01485_),
    .B(_04141_),
    .Y(_04142_)
  );
  NAND _12361_ (
    .A(_01560_),
    .B(_04140_),
    .Y(_04143_)
  );
  NAND _12362_ (
    .A(_04142_),
    .B(_04143_),
    .Y(_04144_)
  );
  OR _12363_ (
    .A(\data_i[2] ),
    .B(_01485_),
    .Y(_04145_)
  );
  AND _12364_ (
    .A(MemWrite_i),
    .B(_04145_),
    .Y(_04146_)
  );
  NAND _12365_ (
    .A(_04144_),
    .B(_04146_),
    .Y(_04147_)
  );
  NAND _12366_ (
    .A(_04134_),
    .B(_04147_),
    .Y(_00146_)
  );
  NAND _12367_ (
    .A(\memory[26][3] ),
    .B(_05361_),
    .Y(_04148_)
  );
  OR _12368_ (
    .A(\memory[26][3] ),
    .B(_01546_),
    .Y(_04149_)
  );
  OR _12369_ (
    .A(\data_i[27] ),
    .B(_01547_),
    .Y(_04150_)
  );
  NAND _12370_ (
    .A(_04149_),
    .B(_04150_),
    .Y(_04151_)
  );
  NAND _12371_ (
    .A(_01551_),
    .B(_04151_),
    .Y(_04152_)
  );
  OR _12372_ (
    .A(\data_i[19] ),
    .B(_01551_),
    .Y(_04153_)
  );
  AND _12373_ (
    .A(_04152_),
    .B(_04153_),
    .Y(_04154_)
  );
  NAND _12374_ (
    .A(\data_i[11] ),
    .B(_01559_),
    .Y(_04155_)
  );
  AND _12375_ (
    .A(_01485_),
    .B(_04155_),
    .Y(_04156_)
  );
  NAND _12376_ (
    .A(_01560_),
    .B(_04154_),
    .Y(_04157_)
  );
  NAND _12377_ (
    .A(_04156_),
    .B(_04157_),
    .Y(_04158_)
  );
  OR _12378_ (
    .A(\data_i[3] ),
    .B(_01485_),
    .Y(_04159_)
  );
  AND _12379_ (
    .A(MemWrite_i),
    .B(_04159_),
    .Y(_04160_)
  );
  NAND _12380_ (
    .A(_04158_),
    .B(_04160_),
    .Y(_04161_)
  );
  NAND _12381_ (
    .A(_04148_),
    .B(_04161_),
    .Y(_00147_)
  );
  NAND _12382_ (
    .A(\memory[26][4] ),
    .B(_05361_),
    .Y(_04162_)
  );
  OR _12383_ (
    .A(\memory[26][4] ),
    .B(_01546_),
    .Y(_04163_)
  );
  OR _12384_ (
    .A(\data_i[28] ),
    .B(_01547_),
    .Y(_04164_)
  );
  NAND _12385_ (
    .A(_04163_),
    .B(_04164_),
    .Y(_04165_)
  );
  NAND _12386_ (
    .A(_01551_),
    .B(_04165_),
    .Y(_04166_)
  );
  OR _12387_ (
    .A(\data_i[20] ),
    .B(_01551_),
    .Y(_04167_)
  );
  AND _12388_ (
    .A(_04166_),
    .B(_04167_),
    .Y(_04168_)
  );
  NAND _12389_ (
    .A(\data_i[12] ),
    .B(_01559_),
    .Y(_04169_)
  );
  AND _12390_ (
    .A(_01485_),
    .B(_04169_),
    .Y(_04170_)
  );
  NAND _12391_ (
    .A(_01560_),
    .B(_04168_),
    .Y(_04171_)
  );
  NAND _12392_ (
    .A(_04170_),
    .B(_04171_),
    .Y(_04172_)
  );
  OR _12393_ (
    .A(\data_i[4] ),
    .B(_01485_),
    .Y(_04173_)
  );
  AND _12394_ (
    .A(MemWrite_i),
    .B(_04173_),
    .Y(_04174_)
  );
  NAND _12395_ (
    .A(_04172_),
    .B(_04174_),
    .Y(_04175_)
  );
  NAND _12396_ (
    .A(_04162_),
    .B(_04175_),
    .Y(_00148_)
  );
  NAND _12397_ (
    .A(\memory[26][5] ),
    .B(_05361_),
    .Y(_04176_)
  );
  OR _12398_ (
    .A(\memory[26][5] ),
    .B(_01546_),
    .Y(_04177_)
  );
  OR _12399_ (
    .A(\data_i[29] ),
    .B(_01547_),
    .Y(_04178_)
  );
  NAND _12400_ (
    .A(_04177_),
    .B(_04178_),
    .Y(_04179_)
  );
  NAND _12401_ (
    .A(_01551_),
    .B(_04179_),
    .Y(_04180_)
  );
  OR _12402_ (
    .A(\data_i[21] ),
    .B(_01551_),
    .Y(_04181_)
  );
  AND _12403_ (
    .A(_04180_),
    .B(_04181_),
    .Y(_04182_)
  );
  NAND _12404_ (
    .A(\data_i[13] ),
    .B(_01559_),
    .Y(_04183_)
  );
  AND _12405_ (
    .A(_01485_),
    .B(_04183_),
    .Y(_04184_)
  );
  NAND _12406_ (
    .A(_01560_),
    .B(_04182_),
    .Y(_04185_)
  );
  NAND _12407_ (
    .A(_04184_),
    .B(_04185_),
    .Y(_04186_)
  );
  OR _12408_ (
    .A(\data_i[5] ),
    .B(_01485_),
    .Y(_04187_)
  );
  AND _12409_ (
    .A(MemWrite_i),
    .B(_04187_),
    .Y(_04188_)
  );
  NAND _12410_ (
    .A(_04186_),
    .B(_04188_),
    .Y(_04189_)
  );
  NAND _12411_ (
    .A(_04176_),
    .B(_04189_),
    .Y(_00149_)
  );
  NAND _12412_ (
    .A(\memory[26][6] ),
    .B(_05361_),
    .Y(_04190_)
  );
  OR _12413_ (
    .A(\memory[26][6] ),
    .B(_01546_),
    .Y(_04191_)
  );
  OR _12414_ (
    .A(\data_i[30] ),
    .B(_01547_),
    .Y(_04192_)
  );
  NAND _12415_ (
    .A(_04191_),
    .B(_04192_),
    .Y(_04193_)
  );
  NAND _12416_ (
    .A(_01551_),
    .B(_04193_),
    .Y(_04194_)
  );
  OR _12417_ (
    .A(\data_i[22] ),
    .B(_01551_),
    .Y(_04195_)
  );
  AND _12418_ (
    .A(_04194_),
    .B(_04195_),
    .Y(_04196_)
  );
  NAND _12419_ (
    .A(\data_i[14] ),
    .B(_01559_),
    .Y(_04197_)
  );
  AND _12420_ (
    .A(_01485_),
    .B(_04197_),
    .Y(_04198_)
  );
  NAND _12421_ (
    .A(_01560_),
    .B(_04196_),
    .Y(_04199_)
  );
  NAND _12422_ (
    .A(_04198_),
    .B(_04199_),
    .Y(_04200_)
  );
  OR _12423_ (
    .A(\data_i[6] ),
    .B(_01485_),
    .Y(_04201_)
  );
  AND _12424_ (
    .A(MemWrite_i),
    .B(_04201_),
    .Y(_04202_)
  );
  NAND _12425_ (
    .A(_04200_),
    .B(_04202_),
    .Y(_04203_)
  );
  NAND _12426_ (
    .A(_04190_),
    .B(_04203_),
    .Y(_00150_)
  );
  NAND _12427_ (
    .A(\memory[26][7] ),
    .B(_05361_),
    .Y(_04204_)
  );
  OR _12428_ (
    .A(\memory[26][7] ),
    .B(_01546_),
    .Y(_04205_)
  );
  OR _12429_ (
    .A(\data_i[31] ),
    .B(_01547_),
    .Y(_04206_)
  );
  NAND _12430_ (
    .A(_04205_),
    .B(_04206_),
    .Y(_04207_)
  );
  NAND _12431_ (
    .A(_01551_),
    .B(_04207_),
    .Y(_04208_)
  );
  OR _12432_ (
    .A(\data_i[23] ),
    .B(_01551_),
    .Y(_04209_)
  );
  AND _12433_ (
    .A(_04208_),
    .B(_04209_),
    .Y(_04210_)
  );
  NAND _12434_ (
    .A(\data_i[15] ),
    .B(_01559_),
    .Y(_04211_)
  );
  AND _12435_ (
    .A(_01485_),
    .B(_04211_),
    .Y(_04212_)
  );
  NAND _12436_ (
    .A(_01560_),
    .B(_04210_),
    .Y(_04213_)
  );
  NAND _12437_ (
    .A(_04212_),
    .B(_04213_),
    .Y(_04214_)
  );
  OR _12438_ (
    .A(\data_i[7] ),
    .B(_01485_),
    .Y(_04215_)
  );
  AND _12439_ (
    .A(MemWrite_i),
    .B(_04215_),
    .Y(_04216_)
  );
  NAND _12440_ (
    .A(_04214_),
    .B(_04216_),
    .Y(_04217_)
  );
  NAND _12441_ (
    .A(_04204_),
    .B(_04217_),
    .Y(_00151_)
  );
  NAND _12442_ (
    .A(\memory[25][0] ),
    .B(_05361_),
    .Y(_04218_)
  );
  OR _12443_ (
    .A(\memory[25][0] ),
    .B(_01469_),
    .Y(_04219_)
  );
  OR _12444_ (
    .A(\data_i[24] ),
    .B(_01470_),
    .Y(_04220_)
  );
  NAND _12445_ (
    .A(_04219_),
    .B(_04220_),
    .Y(_04221_)
  );
  NAND _12446_ (
    .A(_01547_),
    .B(_04221_),
    .Y(_04222_)
  );
  OR _12447_ (
    .A(\data_i[16] ),
    .B(_01547_),
    .Y(_04223_)
  );
  AND _12448_ (
    .A(_04222_),
    .B(_04223_),
    .Y(_04224_)
  );
  NAND _12449_ (
    .A(\data_i[8] ),
    .B(_01550_),
    .Y(_04225_)
  );
  AND _12450_ (
    .A(_01560_),
    .B(_04225_),
    .Y(_04226_)
  );
  NAND _12451_ (
    .A(_01551_),
    .B(_04224_),
    .Y(_04227_)
  );
  NAND _12452_ (
    .A(_04226_),
    .B(_04227_),
    .Y(_04228_)
  );
  OR _12453_ (
    .A(\data_i[0] ),
    .B(_01560_),
    .Y(_04229_)
  );
  AND _12454_ (
    .A(MemWrite_i),
    .B(_04229_),
    .Y(_04230_)
  );
  NAND _12455_ (
    .A(_04228_),
    .B(_04230_),
    .Y(_04231_)
  );
  NAND _12456_ (
    .A(_04218_),
    .B(_04231_),
    .Y(_00136_)
  );
  NAND _12457_ (
    .A(\memory[25][1] ),
    .B(_05361_),
    .Y(_04232_)
  );
  OR _12458_ (
    .A(\memory[25][1] ),
    .B(_01469_),
    .Y(_04233_)
  );
  OR _12459_ (
    .A(\data_i[25] ),
    .B(_01470_),
    .Y(_04234_)
  );
  NAND _12460_ (
    .A(_04233_),
    .B(_04234_),
    .Y(_04235_)
  );
  NAND _12461_ (
    .A(_01547_),
    .B(_04235_),
    .Y(_04236_)
  );
  OR _12462_ (
    .A(\data_i[17] ),
    .B(_01547_),
    .Y(_04237_)
  );
  AND _12463_ (
    .A(_04236_),
    .B(_04237_),
    .Y(_04238_)
  );
  NAND _12464_ (
    .A(\data_i[9] ),
    .B(_01550_),
    .Y(_04239_)
  );
  AND _12465_ (
    .A(_01560_),
    .B(_04239_),
    .Y(_04240_)
  );
  NAND _12466_ (
    .A(_01551_),
    .B(_04238_),
    .Y(_04241_)
  );
  NAND _12467_ (
    .A(_04240_),
    .B(_04241_),
    .Y(_04242_)
  );
  OR _12468_ (
    .A(\data_i[1] ),
    .B(_01560_),
    .Y(_04243_)
  );
  AND _12469_ (
    .A(MemWrite_i),
    .B(_04243_),
    .Y(_04244_)
  );
  NAND _12470_ (
    .A(_04242_),
    .B(_04244_),
    .Y(_04245_)
  );
  NAND _12471_ (
    .A(_04232_),
    .B(_04245_),
    .Y(_00137_)
  );
  NAND _12472_ (
    .A(\memory[25][2] ),
    .B(_05361_),
    .Y(_04246_)
  );
  OR _12473_ (
    .A(\memory[25][2] ),
    .B(_01469_),
    .Y(_04247_)
  );
  OR _12474_ (
    .A(\data_i[26] ),
    .B(_01470_),
    .Y(_04248_)
  );
  NAND _12475_ (
    .A(_04247_),
    .B(_04248_),
    .Y(_04249_)
  );
  NAND _12476_ (
    .A(_01547_),
    .B(_04249_),
    .Y(_04250_)
  );
  OR _12477_ (
    .A(\data_i[18] ),
    .B(_01547_),
    .Y(_04251_)
  );
  AND _12478_ (
    .A(_04250_),
    .B(_04251_),
    .Y(_04252_)
  );
  NAND _12479_ (
    .A(\data_i[10] ),
    .B(_01550_),
    .Y(_04253_)
  );
  AND _12480_ (
    .A(_01560_),
    .B(_04253_),
    .Y(_04254_)
  );
  NAND _12481_ (
    .A(_01551_),
    .B(_04252_),
    .Y(_04255_)
  );
  NAND _12482_ (
    .A(_04254_),
    .B(_04255_),
    .Y(_04256_)
  );
  OR _12483_ (
    .A(\data_i[2] ),
    .B(_01560_),
    .Y(_04257_)
  );
  AND _12484_ (
    .A(MemWrite_i),
    .B(_04257_),
    .Y(_04258_)
  );
  NAND _12485_ (
    .A(_04256_),
    .B(_04258_),
    .Y(_04259_)
  );
  NAND _12486_ (
    .A(_04246_),
    .B(_04259_),
    .Y(_00138_)
  );
  NAND _12487_ (
    .A(\memory[25][3] ),
    .B(_05361_),
    .Y(_04260_)
  );
  OR _12488_ (
    .A(\memory[25][3] ),
    .B(_01469_),
    .Y(_04261_)
  );
  OR _12489_ (
    .A(\data_i[27] ),
    .B(_01470_),
    .Y(_04262_)
  );
  NAND _12490_ (
    .A(_04261_),
    .B(_04262_),
    .Y(_04263_)
  );
  NAND _12491_ (
    .A(_01547_),
    .B(_04263_),
    .Y(_04264_)
  );
  OR _12492_ (
    .A(\data_i[19] ),
    .B(_01547_),
    .Y(_04265_)
  );
  AND _12493_ (
    .A(_04264_),
    .B(_04265_),
    .Y(_04266_)
  );
  NAND _12494_ (
    .A(\data_i[11] ),
    .B(_01550_),
    .Y(_04267_)
  );
  AND _12495_ (
    .A(_01560_),
    .B(_04267_),
    .Y(_04268_)
  );
  NAND _12496_ (
    .A(_01551_),
    .B(_04266_),
    .Y(_04269_)
  );
  NAND _12497_ (
    .A(_04268_),
    .B(_04269_),
    .Y(_04270_)
  );
  OR _12498_ (
    .A(\data_i[3] ),
    .B(_01560_),
    .Y(_04271_)
  );
  AND _12499_ (
    .A(MemWrite_i),
    .B(_04271_),
    .Y(_04272_)
  );
  NAND _12500_ (
    .A(_04270_),
    .B(_04272_),
    .Y(_04273_)
  );
  NAND _12501_ (
    .A(_04260_),
    .B(_04273_),
    .Y(_00139_)
  );
  NAND _12502_ (
    .A(\memory[25][4] ),
    .B(_05361_),
    .Y(_04274_)
  );
  OR _12503_ (
    .A(\memory[25][4] ),
    .B(_01469_),
    .Y(_04275_)
  );
  OR _12504_ (
    .A(\data_i[28] ),
    .B(_01470_),
    .Y(_04276_)
  );
  NAND _12505_ (
    .A(_04275_),
    .B(_04276_),
    .Y(_04277_)
  );
  NAND _12506_ (
    .A(_01547_),
    .B(_04277_),
    .Y(_04278_)
  );
  OR _12507_ (
    .A(\data_i[20] ),
    .B(_01547_),
    .Y(_04279_)
  );
  AND _12508_ (
    .A(_04278_),
    .B(_04279_),
    .Y(_04280_)
  );
  NAND _12509_ (
    .A(\data_i[12] ),
    .B(_01550_),
    .Y(_04281_)
  );
  AND _12510_ (
    .A(_01560_),
    .B(_04281_),
    .Y(_04282_)
  );
  NAND _12511_ (
    .A(_01551_),
    .B(_04280_),
    .Y(_04283_)
  );
  NAND _12512_ (
    .A(_04282_),
    .B(_04283_),
    .Y(_04284_)
  );
  OR _12513_ (
    .A(\data_i[4] ),
    .B(_01560_),
    .Y(_04285_)
  );
  AND _12514_ (
    .A(MemWrite_i),
    .B(_04285_),
    .Y(_04286_)
  );
  NAND _12515_ (
    .A(_04284_),
    .B(_04286_),
    .Y(_04287_)
  );
  NAND _12516_ (
    .A(_04274_),
    .B(_04287_),
    .Y(_00140_)
  );
  NAND _12517_ (
    .A(\memory[25][5] ),
    .B(_05361_),
    .Y(_04288_)
  );
  OR _12518_ (
    .A(\memory[25][5] ),
    .B(_01469_),
    .Y(_04289_)
  );
  OR _12519_ (
    .A(\data_i[29] ),
    .B(_01470_),
    .Y(_04290_)
  );
  NAND _12520_ (
    .A(_04289_),
    .B(_04290_),
    .Y(_04291_)
  );
  NAND _12521_ (
    .A(_01547_),
    .B(_04291_),
    .Y(_04292_)
  );
  OR _12522_ (
    .A(\data_i[21] ),
    .B(_01547_),
    .Y(_04293_)
  );
  AND _12523_ (
    .A(_04292_),
    .B(_04293_),
    .Y(_04294_)
  );
  NAND _12524_ (
    .A(\data_i[13] ),
    .B(_01550_),
    .Y(_04295_)
  );
  AND _12525_ (
    .A(_01560_),
    .B(_04295_),
    .Y(_04296_)
  );
  NAND _12526_ (
    .A(_01551_),
    .B(_04294_),
    .Y(_04297_)
  );
  NAND _12527_ (
    .A(_04296_),
    .B(_04297_),
    .Y(_04298_)
  );
  OR _12528_ (
    .A(\data_i[5] ),
    .B(_01560_),
    .Y(_04299_)
  );
  AND _12529_ (
    .A(MemWrite_i),
    .B(_04299_),
    .Y(_04300_)
  );
  NAND _12530_ (
    .A(_04298_),
    .B(_04300_),
    .Y(_04301_)
  );
  NAND _12531_ (
    .A(_04288_),
    .B(_04301_),
    .Y(_00141_)
  );
  NAND _12532_ (
    .A(\memory[25][6] ),
    .B(_05361_),
    .Y(_04302_)
  );
  OR _12533_ (
    .A(\memory[25][6] ),
    .B(_01469_),
    .Y(_04303_)
  );
  OR _12534_ (
    .A(\data_i[30] ),
    .B(_01470_),
    .Y(_04304_)
  );
  NAND _12535_ (
    .A(_04303_),
    .B(_04304_),
    .Y(_04305_)
  );
  NAND _12536_ (
    .A(_01547_),
    .B(_04305_),
    .Y(_04306_)
  );
  OR _12537_ (
    .A(\data_i[22] ),
    .B(_01547_),
    .Y(_04307_)
  );
  AND _12538_ (
    .A(_04306_),
    .B(_04307_),
    .Y(_04308_)
  );
  NAND _12539_ (
    .A(\data_i[14] ),
    .B(_01550_),
    .Y(_04309_)
  );
  AND _12540_ (
    .A(_01560_),
    .B(_04309_),
    .Y(_04310_)
  );
  NAND _12541_ (
    .A(_01551_),
    .B(_04308_),
    .Y(_04311_)
  );
  NAND _12542_ (
    .A(_04310_),
    .B(_04311_),
    .Y(_04312_)
  );
  OR _12543_ (
    .A(\data_i[6] ),
    .B(_01560_),
    .Y(_04313_)
  );
  AND _12544_ (
    .A(MemWrite_i),
    .B(_04313_),
    .Y(_04314_)
  );
  NAND _12545_ (
    .A(_04312_),
    .B(_04314_),
    .Y(_04315_)
  );
  NAND _12546_ (
    .A(_04302_),
    .B(_04315_),
    .Y(_00142_)
  );
  NAND _12547_ (
    .A(\memory[25][7] ),
    .B(_05361_),
    .Y(_04316_)
  );
  OR _12548_ (
    .A(\memory[25][7] ),
    .B(_01469_),
    .Y(_04317_)
  );
  OR _12549_ (
    .A(\data_i[31] ),
    .B(_01470_),
    .Y(_04318_)
  );
  NAND _12550_ (
    .A(_04317_),
    .B(_04318_),
    .Y(_04319_)
  );
  NAND _12551_ (
    .A(_01547_),
    .B(_04319_),
    .Y(_04320_)
  );
  OR _12552_ (
    .A(\data_i[23] ),
    .B(_01547_),
    .Y(_04321_)
  );
  AND _12553_ (
    .A(_04320_),
    .B(_04321_),
    .Y(_04322_)
  );
  NAND _12554_ (
    .A(\data_i[15] ),
    .B(_01550_),
    .Y(_04323_)
  );
  AND _12555_ (
    .A(_01560_),
    .B(_04323_),
    .Y(_04324_)
  );
  NAND _12556_ (
    .A(_01551_),
    .B(_04322_),
    .Y(_04325_)
  );
  NAND _12557_ (
    .A(_04324_),
    .B(_04325_),
    .Y(_04326_)
  );
  OR _12558_ (
    .A(\data_i[7] ),
    .B(_01560_),
    .Y(_04327_)
  );
  AND _12559_ (
    .A(MemWrite_i),
    .B(_04327_),
    .Y(_04328_)
  );
  NAND _12560_ (
    .A(_04326_),
    .B(_04328_),
    .Y(_04329_)
  );
  NAND _12561_ (
    .A(_04316_),
    .B(_04329_),
    .Y(_00143_)
  );
  NAND _12562_ (
    .A(\memory[24][0] ),
    .B(_05361_),
    .Y(_04330_)
  );
  OR _12563_ (
    .A(\memory[24][0] ),
    .B(_01474_),
    .Y(_04331_)
  );
  OR _12564_ (
    .A(\data_i[24] ),
    .B(_01475_),
    .Y(_04332_)
  );
  NAND _12565_ (
    .A(_04331_),
    .B(_04332_),
    .Y(_04333_)
  );
  NAND _12566_ (
    .A(_01470_),
    .B(_04333_),
    .Y(_04334_)
  );
  OR _12567_ (
    .A(\data_i[16] ),
    .B(_01470_),
    .Y(_04335_)
  );
  AND _12568_ (
    .A(_04334_),
    .B(_04335_),
    .Y(_04336_)
  );
  NAND _12569_ (
    .A(\data_i[8] ),
    .B(_01546_),
    .Y(_04337_)
  );
  AND _12570_ (
    .A(_01551_),
    .B(_04337_),
    .Y(_04338_)
  );
  NAND _12571_ (
    .A(_01547_),
    .B(_04336_),
    .Y(_04339_)
  );
  NAND _12572_ (
    .A(_04338_),
    .B(_04339_),
    .Y(_04340_)
  );
  OR _12573_ (
    .A(\data_i[0] ),
    .B(_01551_),
    .Y(_04341_)
  );
  AND _12574_ (
    .A(MemWrite_i),
    .B(_04341_),
    .Y(_04342_)
  );
  NAND _12575_ (
    .A(_04340_),
    .B(_04342_),
    .Y(_04343_)
  );
  NAND _12576_ (
    .A(_04330_),
    .B(_04343_),
    .Y(_00128_)
  );
  NAND _12577_ (
    .A(\memory[24][1] ),
    .B(_05361_),
    .Y(_04344_)
  );
  OR _12578_ (
    .A(\memory[24][1] ),
    .B(_01474_),
    .Y(_04345_)
  );
  OR _12579_ (
    .A(\data_i[25] ),
    .B(_01475_),
    .Y(_04346_)
  );
  NAND _12580_ (
    .A(_04345_),
    .B(_04346_),
    .Y(_04347_)
  );
  NAND _12581_ (
    .A(_01470_),
    .B(_04347_),
    .Y(_04348_)
  );
  OR _12582_ (
    .A(\data_i[17] ),
    .B(_01470_),
    .Y(_04349_)
  );
  AND _12583_ (
    .A(_04348_),
    .B(_04349_),
    .Y(_04350_)
  );
  NAND _12584_ (
    .A(\data_i[9] ),
    .B(_01546_),
    .Y(_04351_)
  );
  AND _12585_ (
    .A(_01551_),
    .B(_04351_),
    .Y(_04352_)
  );
  NAND _12586_ (
    .A(_01547_),
    .B(_04350_),
    .Y(_04353_)
  );
  NAND _12587_ (
    .A(_04352_),
    .B(_04353_),
    .Y(_04354_)
  );
  OR _12588_ (
    .A(\data_i[1] ),
    .B(_01551_),
    .Y(_04355_)
  );
  AND _12589_ (
    .A(MemWrite_i),
    .B(_04355_),
    .Y(_04356_)
  );
  NAND _12590_ (
    .A(_04354_),
    .B(_04356_),
    .Y(_04357_)
  );
  NAND _12591_ (
    .A(_04344_),
    .B(_04357_),
    .Y(_00129_)
  );
  NAND _12592_ (
    .A(\memory[24][2] ),
    .B(_05361_),
    .Y(_04358_)
  );
  OR _12593_ (
    .A(\memory[24][2] ),
    .B(_01474_),
    .Y(_04359_)
  );
  OR _12594_ (
    .A(\data_i[26] ),
    .B(_01475_),
    .Y(_04360_)
  );
  NAND _12595_ (
    .A(_04359_),
    .B(_04360_),
    .Y(_04361_)
  );
  NAND _12596_ (
    .A(_01470_),
    .B(_04361_),
    .Y(_04362_)
  );
  OR _12597_ (
    .A(\data_i[18] ),
    .B(_01470_),
    .Y(_04363_)
  );
  AND _12598_ (
    .A(_04362_),
    .B(_04363_),
    .Y(_04364_)
  );
  NAND _12599_ (
    .A(\data_i[10] ),
    .B(_01546_),
    .Y(_04365_)
  );
  AND _12600_ (
    .A(_01551_),
    .B(_04365_),
    .Y(_04366_)
  );
  NAND _12601_ (
    .A(_01547_),
    .B(_04364_),
    .Y(_04367_)
  );
  NAND _12602_ (
    .A(_04366_),
    .B(_04367_),
    .Y(_04368_)
  );
  OR _12603_ (
    .A(\data_i[2] ),
    .B(_01551_),
    .Y(_04369_)
  );
  AND _12604_ (
    .A(MemWrite_i),
    .B(_04369_),
    .Y(_04370_)
  );
  NAND _12605_ (
    .A(_04368_),
    .B(_04370_),
    .Y(_04371_)
  );
  NAND _12606_ (
    .A(_04358_),
    .B(_04371_),
    .Y(_00130_)
  );
  NAND _12607_ (
    .A(\memory[24][3] ),
    .B(_05361_),
    .Y(_04372_)
  );
  OR _12608_ (
    .A(\memory[24][3] ),
    .B(_01474_),
    .Y(_04373_)
  );
  OR _12609_ (
    .A(\data_i[27] ),
    .B(_01475_),
    .Y(_04374_)
  );
  NAND _12610_ (
    .A(_04373_),
    .B(_04374_),
    .Y(_04375_)
  );
  NAND _12611_ (
    .A(_01470_),
    .B(_04375_),
    .Y(_04376_)
  );
  OR _12612_ (
    .A(\data_i[19] ),
    .B(_01470_),
    .Y(_04377_)
  );
  AND _12613_ (
    .A(_04376_),
    .B(_04377_),
    .Y(_04378_)
  );
  NAND _12614_ (
    .A(\data_i[11] ),
    .B(_01546_),
    .Y(_04379_)
  );
  AND _12615_ (
    .A(_01551_),
    .B(_04379_),
    .Y(_04380_)
  );
  NAND _12616_ (
    .A(_01547_),
    .B(_04378_),
    .Y(_04381_)
  );
  NAND _12617_ (
    .A(_04380_),
    .B(_04381_),
    .Y(_04382_)
  );
  OR _12618_ (
    .A(\data_i[3] ),
    .B(_01551_),
    .Y(_04383_)
  );
  AND _12619_ (
    .A(MemWrite_i),
    .B(_04383_),
    .Y(_04384_)
  );
  NAND _12620_ (
    .A(_04382_),
    .B(_04384_),
    .Y(_04385_)
  );
  NAND _12621_ (
    .A(_04372_),
    .B(_04385_),
    .Y(_00131_)
  );
  NAND _12622_ (
    .A(\memory[24][4] ),
    .B(_05361_),
    .Y(_04386_)
  );
  OR _12623_ (
    .A(\memory[24][4] ),
    .B(_01474_),
    .Y(_04387_)
  );
  OR _12624_ (
    .A(\data_i[28] ),
    .B(_01475_),
    .Y(_04388_)
  );
  NAND _12625_ (
    .A(_04387_),
    .B(_04388_),
    .Y(_04389_)
  );
  NAND _12626_ (
    .A(_01470_),
    .B(_04389_),
    .Y(_04390_)
  );
  OR _12627_ (
    .A(\data_i[20] ),
    .B(_01470_),
    .Y(_04391_)
  );
  AND _12628_ (
    .A(_04390_),
    .B(_04391_),
    .Y(_04392_)
  );
  NAND _12629_ (
    .A(\data_i[12] ),
    .B(_01546_),
    .Y(_04393_)
  );
  AND _12630_ (
    .A(_01551_),
    .B(_04393_),
    .Y(_04394_)
  );
  NAND _12631_ (
    .A(_01547_),
    .B(_04392_),
    .Y(_04395_)
  );
  NAND _12632_ (
    .A(_04394_),
    .B(_04395_),
    .Y(_04396_)
  );
  OR _12633_ (
    .A(\data_i[4] ),
    .B(_01551_),
    .Y(_04397_)
  );
  AND _12634_ (
    .A(MemWrite_i),
    .B(_04397_),
    .Y(_04398_)
  );
  NAND _12635_ (
    .A(_04396_),
    .B(_04398_),
    .Y(_04399_)
  );
  NAND _12636_ (
    .A(_04386_),
    .B(_04399_),
    .Y(_00132_)
  );
  NAND _12637_ (
    .A(\memory[24][5] ),
    .B(_05361_),
    .Y(_04400_)
  );
  OR _12638_ (
    .A(\memory[24][5] ),
    .B(_01474_),
    .Y(_04401_)
  );
  OR _12639_ (
    .A(\data_i[29] ),
    .B(_01475_),
    .Y(_04402_)
  );
  NAND _12640_ (
    .A(_04401_),
    .B(_04402_),
    .Y(_04403_)
  );
  NAND _12641_ (
    .A(_01470_),
    .B(_04403_),
    .Y(_04404_)
  );
  OR _12642_ (
    .A(\data_i[21] ),
    .B(_01470_),
    .Y(_04405_)
  );
  AND _12643_ (
    .A(_04404_),
    .B(_04405_),
    .Y(_04406_)
  );
  NAND _12644_ (
    .A(\data_i[13] ),
    .B(_01546_),
    .Y(_04407_)
  );
  AND _12645_ (
    .A(_01551_),
    .B(_04407_),
    .Y(_04408_)
  );
  NAND _12646_ (
    .A(_01547_),
    .B(_04406_),
    .Y(_04409_)
  );
  NAND _12647_ (
    .A(_04408_),
    .B(_04409_),
    .Y(_04410_)
  );
  OR _12648_ (
    .A(\data_i[5] ),
    .B(_01551_),
    .Y(_04411_)
  );
  AND _12649_ (
    .A(MemWrite_i),
    .B(_04411_),
    .Y(_04412_)
  );
  NAND _12650_ (
    .A(_04410_),
    .B(_04412_),
    .Y(_04413_)
  );
  NAND _12651_ (
    .A(_04400_),
    .B(_04413_),
    .Y(_00133_)
  );
  NAND _12652_ (
    .A(\memory[24][6] ),
    .B(_05361_),
    .Y(_04414_)
  );
  OR _12653_ (
    .A(\memory[24][6] ),
    .B(_01474_),
    .Y(_04415_)
  );
  OR _12654_ (
    .A(\data_i[30] ),
    .B(_01475_),
    .Y(_04416_)
  );
  NAND _12655_ (
    .A(_04415_),
    .B(_04416_),
    .Y(_04417_)
  );
  NAND _12656_ (
    .A(_01470_),
    .B(_04417_),
    .Y(_04418_)
  );
  OR _12657_ (
    .A(\data_i[22] ),
    .B(_01470_),
    .Y(_04419_)
  );
  AND _12658_ (
    .A(_04418_),
    .B(_04419_),
    .Y(_04420_)
  );
  NAND _12659_ (
    .A(\data_i[14] ),
    .B(_01546_),
    .Y(_04421_)
  );
  AND _12660_ (
    .A(_01551_),
    .B(_04421_),
    .Y(_04422_)
  );
  NAND _12661_ (
    .A(_01547_),
    .B(_04420_),
    .Y(_04423_)
  );
  NAND _12662_ (
    .A(_04422_),
    .B(_04423_),
    .Y(_04424_)
  );
  OR _12663_ (
    .A(\data_i[6] ),
    .B(_01551_),
    .Y(_04425_)
  );
  AND _12664_ (
    .A(MemWrite_i),
    .B(_04425_),
    .Y(_04426_)
  );
  NAND _12665_ (
    .A(_04424_),
    .B(_04426_),
    .Y(_04427_)
  );
  NAND _12666_ (
    .A(_04414_),
    .B(_04427_),
    .Y(_00134_)
  );
  NAND _12667_ (
    .A(\memory[24][7] ),
    .B(_05361_),
    .Y(_04428_)
  );
  OR _12668_ (
    .A(\memory[24][7] ),
    .B(_01474_),
    .Y(_04429_)
  );
  OR _12669_ (
    .A(\data_i[31] ),
    .B(_01475_),
    .Y(_04430_)
  );
  NAND _12670_ (
    .A(_04429_),
    .B(_04430_),
    .Y(_04431_)
  );
  NAND _12671_ (
    .A(_01470_),
    .B(_04431_),
    .Y(_04432_)
  );
  OR _12672_ (
    .A(\data_i[23] ),
    .B(_01470_),
    .Y(_04433_)
  );
  AND _12673_ (
    .A(_04432_),
    .B(_04433_),
    .Y(_04434_)
  );
  NAND _12674_ (
    .A(\data_i[15] ),
    .B(_01546_),
    .Y(_04435_)
  );
  AND _12675_ (
    .A(_01551_),
    .B(_04435_),
    .Y(_04436_)
  );
  NAND _12676_ (
    .A(_01547_),
    .B(_04434_),
    .Y(_04437_)
  );
  NAND _12677_ (
    .A(_04436_),
    .B(_04437_),
    .Y(_04438_)
  );
  OR _12678_ (
    .A(\data_i[7] ),
    .B(_01551_),
    .Y(_04439_)
  );
  AND _12679_ (
    .A(MemWrite_i),
    .B(_04439_),
    .Y(_04440_)
  );
  NAND _12680_ (
    .A(_04438_),
    .B(_04440_),
    .Y(_04441_)
  );
  NAND _12681_ (
    .A(_04428_),
    .B(_04441_),
    .Y(_00135_)
  );
  NAND _12682_ (
    .A(\memory[23][0] ),
    .B(_05361_),
    .Y(_04442_)
  );
  OR _12683_ (
    .A(\memory[23][0] ),
    .B(_01553_),
    .Y(_04443_)
  );
  OR _12684_ (
    .A(\data_i[24] ),
    .B(_01554_),
    .Y(_04444_)
  );
  NAND _12685_ (
    .A(_04443_),
    .B(_04444_),
    .Y(_04445_)
  );
  NAND _12686_ (
    .A(_01475_),
    .B(_04445_),
    .Y(_04446_)
  );
  OR _12687_ (
    .A(\data_i[16] ),
    .B(_01475_),
    .Y(_04447_)
  );
  AND _12688_ (
    .A(_04446_),
    .B(_04447_),
    .Y(_04448_)
  );
  NAND _12689_ (
    .A(\data_i[8] ),
    .B(_01469_),
    .Y(_04449_)
  );
  AND _12690_ (
    .A(_01547_),
    .B(_04449_),
    .Y(_04450_)
  );
  NAND _12691_ (
    .A(_01470_),
    .B(_04448_),
    .Y(_04451_)
  );
  NAND _12692_ (
    .A(_04450_),
    .B(_04451_),
    .Y(_04452_)
  );
  OR _12693_ (
    .A(\data_i[0] ),
    .B(_01547_),
    .Y(_04453_)
  );
  AND _12694_ (
    .A(MemWrite_i),
    .B(_04453_),
    .Y(_04454_)
  );
  NAND _12695_ (
    .A(_04452_),
    .B(_04454_),
    .Y(_04455_)
  );
  NAND _12696_ (
    .A(_04442_),
    .B(_04455_),
    .Y(_00120_)
  );
  NAND _12697_ (
    .A(\memory[23][1] ),
    .B(_05361_),
    .Y(_04456_)
  );
  OR _12698_ (
    .A(\memory[23][1] ),
    .B(_01553_),
    .Y(_04457_)
  );
  OR _12699_ (
    .A(\data_i[25] ),
    .B(_01554_),
    .Y(_04458_)
  );
  NAND _12700_ (
    .A(_04457_),
    .B(_04458_),
    .Y(_04459_)
  );
  NAND _12701_ (
    .A(_01475_),
    .B(_04459_),
    .Y(_04460_)
  );
  OR _12702_ (
    .A(\data_i[17] ),
    .B(_01475_),
    .Y(_04461_)
  );
  AND _12703_ (
    .A(_04460_),
    .B(_04461_),
    .Y(_04462_)
  );
  NAND _12704_ (
    .A(\data_i[9] ),
    .B(_01469_),
    .Y(_04463_)
  );
  AND _12705_ (
    .A(_01547_),
    .B(_04463_),
    .Y(_04464_)
  );
  NAND _12706_ (
    .A(_01470_),
    .B(_04462_),
    .Y(_04465_)
  );
  NAND _12707_ (
    .A(_04464_),
    .B(_04465_),
    .Y(_04466_)
  );
  OR _12708_ (
    .A(\data_i[1] ),
    .B(_01547_),
    .Y(_04467_)
  );
  AND _12709_ (
    .A(MemWrite_i),
    .B(_04467_),
    .Y(_04468_)
  );
  NAND _12710_ (
    .A(_04466_),
    .B(_04468_),
    .Y(_04469_)
  );
  NAND _12711_ (
    .A(_04456_),
    .B(_04469_),
    .Y(_00121_)
  );
  NAND _12712_ (
    .A(\memory[23][2] ),
    .B(_05361_),
    .Y(_04470_)
  );
  OR _12713_ (
    .A(\memory[23][2] ),
    .B(_01553_),
    .Y(_04471_)
  );
  OR _12714_ (
    .A(\data_i[26] ),
    .B(_01554_),
    .Y(_04472_)
  );
  NAND _12715_ (
    .A(_04471_),
    .B(_04472_),
    .Y(_04473_)
  );
  NAND _12716_ (
    .A(_01475_),
    .B(_04473_),
    .Y(_04474_)
  );
  OR _12717_ (
    .A(\data_i[18] ),
    .B(_01475_),
    .Y(_04475_)
  );
  AND _12718_ (
    .A(_04474_),
    .B(_04475_),
    .Y(_04476_)
  );
  NAND _12719_ (
    .A(\data_i[10] ),
    .B(_01469_),
    .Y(_04477_)
  );
  AND _12720_ (
    .A(_01547_),
    .B(_04477_),
    .Y(_04478_)
  );
  NAND _12721_ (
    .A(_01470_),
    .B(_04476_),
    .Y(_04479_)
  );
  NAND _12722_ (
    .A(_04478_),
    .B(_04479_),
    .Y(_04480_)
  );
  OR _12723_ (
    .A(\data_i[2] ),
    .B(_01547_),
    .Y(_04481_)
  );
  AND _12724_ (
    .A(MemWrite_i),
    .B(_04481_),
    .Y(_04482_)
  );
  NAND _12725_ (
    .A(_04480_),
    .B(_04482_),
    .Y(_04483_)
  );
  NAND _12726_ (
    .A(_04470_),
    .B(_04483_),
    .Y(_00122_)
  );
  NAND _12727_ (
    .A(\memory[23][3] ),
    .B(_05361_),
    .Y(_04484_)
  );
  OR _12728_ (
    .A(\memory[23][3] ),
    .B(_01553_),
    .Y(_04485_)
  );
  OR _12729_ (
    .A(\data_i[27] ),
    .B(_01554_),
    .Y(_04486_)
  );
  NAND _12730_ (
    .A(_04485_),
    .B(_04486_),
    .Y(_04487_)
  );
  NAND _12731_ (
    .A(_01475_),
    .B(_04487_),
    .Y(_04488_)
  );
  OR _12732_ (
    .A(\data_i[19] ),
    .B(_01475_),
    .Y(_04489_)
  );
  AND _12733_ (
    .A(_04488_),
    .B(_04489_),
    .Y(_04490_)
  );
  NAND _12734_ (
    .A(\data_i[11] ),
    .B(_01469_),
    .Y(_04491_)
  );
  AND _12735_ (
    .A(_01547_),
    .B(_04491_),
    .Y(_04492_)
  );
  NAND _12736_ (
    .A(_01470_),
    .B(_04490_),
    .Y(_04493_)
  );
  NAND _12737_ (
    .A(_04492_),
    .B(_04493_),
    .Y(_04494_)
  );
  OR _12738_ (
    .A(\data_i[3] ),
    .B(_01547_),
    .Y(_04495_)
  );
  AND _12739_ (
    .A(MemWrite_i),
    .B(_04495_),
    .Y(_04496_)
  );
  NAND _12740_ (
    .A(_04494_),
    .B(_04496_),
    .Y(_04497_)
  );
  NAND _12741_ (
    .A(_04484_),
    .B(_04497_),
    .Y(_00123_)
  );
  NAND _12742_ (
    .A(\memory[23][4] ),
    .B(_05361_),
    .Y(_04498_)
  );
  OR _12743_ (
    .A(\memory[23][4] ),
    .B(_01553_),
    .Y(_04499_)
  );
  OR _12744_ (
    .A(\data_i[28] ),
    .B(_01554_),
    .Y(_04500_)
  );
  NAND _12745_ (
    .A(_04499_),
    .B(_04500_),
    .Y(_04501_)
  );
  NAND _12746_ (
    .A(_01475_),
    .B(_04501_),
    .Y(_04502_)
  );
  OR _12747_ (
    .A(\data_i[20] ),
    .B(_01475_),
    .Y(_04503_)
  );
  AND _12748_ (
    .A(_04502_),
    .B(_04503_),
    .Y(_04504_)
  );
  NAND _12749_ (
    .A(\data_i[12] ),
    .B(_01469_),
    .Y(_04505_)
  );
  AND _12750_ (
    .A(_01547_),
    .B(_04505_),
    .Y(_04506_)
  );
  NAND _12751_ (
    .A(_01470_),
    .B(_04504_),
    .Y(_04507_)
  );
  NAND _12752_ (
    .A(_04506_),
    .B(_04507_),
    .Y(_04508_)
  );
  OR _12753_ (
    .A(\data_i[4] ),
    .B(_01547_),
    .Y(_04509_)
  );
  AND _12754_ (
    .A(MemWrite_i),
    .B(_04509_),
    .Y(_04510_)
  );
  NAND _12755_ (
    .A(_04508_),
    .B(_04510_),
    .Y(_04511_)
  );
  NAND _12756_ (
    .A(_04498_),
    .B(_04511_),
    .Y(_00124_)
  );
  NAND _12757_ (
    .A(\memory[23][5] ),
    .B(_05361_),
    .Y(_04512_)
  );
  OR _12758_ (
    .A(\memory[23][5] ),
    .B(_01553_),
    .Y(_04513_)
  );
  OR _12759_ (
    .A(\data_i[29] ),
    .B(_01554_),
    .Y(_04514_)
  );
  NAND _12760_ (
    .A(_04513_),
    .B(_04514_),
    .Y(_04515_)
  );
  NAND _12761_ (
    .A(_01475_),
    .B(_04515_),
    .Y(_04516_)
  );
  OR _12762_ (
    .A(\data_i[21] ),
    .B(_01475_),
    .Y(_04517_)
  );
  AND _12763_ (
    .A(_04516_),
    .B(_04517_),
    .Y(_04518_)
  );
  NAND _12764_ (
    .A(\data_i[13] ),
    .B(_01469_),
    .Y(_04519_)
  );
  AND _12765_ (
    .A(_01547_),
    .B(_04519_),
    .Y(_04520_)
  );
  NAND _12766_ (
    .A(_01470_),
    .B(_04518_),
    .Y(_04521_)
  );
  NAND _12767_ (
    .A(_04520_),
    .B(_04521_),
    .Y(_04522_)
  );
  OR _12768_ (
    .A(\data_i[5] ),
    .B(_01547_),
    .Y(_04523_)
  );
  AND _12769_ (
    .A(MemWrite_i),
    .B(_04523_),
    .Y(_04524_)
  );
  NAND _12770_ (
    .A(_04522_),
    .B(_04524_),
    .Y(_04525_)
  );
  NAND _12771_ (
    .A(_04512_),
    .B(_04525_),
    .Y(_00125_)
  );
  NAND _12772_ (
    .A(\memory[23][6] ),
    .B(_05361_),
    .Y(_04526_)
  );
  OR _12773_ (
    .A(\memory[23][6] ),
    .B(_01553_),
    .Y(_04527_)
  );
  OR _12774_ (
    .A(\data_i[30] ),
    .B(_01554_),
    .Y(_04528_)
  );
  NAND _12775_ (
    .A(_04527_),
    .B(_04528_),
    .Y(_04529_)
  );
  NAND _12776_ (
    .A(_01475_),
    .B(_04529_),
    .Y(_04530_)
  );
  OR _12777_ (
    .A(\data_i[22] ),
    .B(_01475_),
    .Y(_04531_)
  );
  AND _12778_ (
    .A(_04530_),
    .B(_04531_),
    .Y(_04532_)
  );
  NAND _12779_ (
    .A(\data_i[14] ),
    .B(_01469_),
    .Y(_04533_)
  );
  AND _12780_ (
    .A(_01547_),
    .B(_04533_),
    .Y(_04534_)
  );
  NAND _12781_ (
    .A(_01470_),
    .B(_04532_),
    .Y(_04535_)
  );
  NAND _12782_ (
    .A(_04534_),
    .B(_04535_),
    .Y(_04536_)
  );
  OR _12783_ (
    .A(\data_i[6] ),
    .B(_01547_),
    .Y(_04537_)
  );
  AND _12784_ (
    .A(MemWrite_i),
    .B(_04537_),
    .Y(_04538_)
  );
  NAND _12785_ (
    .A(_04536_),
    .B(_04538_),
    .Y(_04539_)
  );
  NAND _12786_ (
    .A(_04526_),
    .B(_04539_),
    .Y(_00126_)
  );
  NAND _12787_ (
    .A(\memory[23][7] ),
    .B(_05361_),
    .Y(_04540_)
  );
  OR _12788_ (
    .A(\memory[23][7] ),
    .B(_01553_),
    .Y(_04541_)
  );
  OR _12789_ (
    .A(\data_i[31] ),
    .B(_01554_),
    .Y(_04542_)
  );
  NAND _12790_ (
    .A(_04541_),
    .B(_04542_),
    .Y(_04543_)
  );
  NAND _12791_ (
    .A(_01475_),
    .B(_04543_),
    .Y(_04544_)
  );
  OR _12792_ (
    .A(\data_i[23] ),
    .B(_01475_),
    .Y(_04545_)
  );
  AND _12793_ (
    .A(_04544_),
    .B(_04545_),
    .Y(_04546_)
  );
  NAND _12794_ (
    .A(\data_i[15] ),
    .B(_01469_),
    .Y(_04547_)
  );
  AND _12795_ (
    .A(_01547_),
    .B(_04547_),
    .Y(_04548_)
  );
  NAND _12796_ (
    .A(_01470_),
    .B(_04546_),
    .Y(_04549_)
  );
  NAND _12797_ (
    .A(_04548_),
    .B(_04549_),
    .Y(_04550_)
  );
  OR _12798_ (
    .A(\data_i[7] ),
    .B(_01547_),
    .Y(_04551_)
  );
  AND _12799_ (
    .A(MemWrite_i),
    .B(_04551_),
    .Y(_04552_)
  );
  NAND _12800_ (
    .A(_04550_),
    .B(_04552_),
    .Y(_04553_)
  );
  NAND _12801_ (
    .A(_04540_),
    .B(_04553_),
    .Y(_00127_)
  );
  NAND _12802_ (
    .A(\memory[22][0] ),
    .B(_05361_),
    .Y(_04554_)
  );
  OR _12803_ (
    .A(\memory[22][0] ),
    .B(_01534_),
    .Y(_04555_)
  );
  OR _12804_ (
    .A(\data_i[24] ),
    .B(_01535_),
    .Y(_04556_)
  );
  NAND _12805_ (
    .A(_04555_),
    .B(_04556_),
    .Y(_04557_)
  );
  NAND _12806_ (
    .A(_01554_),
    .B(_04557_),
    .Y(_04558_)
  );
  OR _12807_ (
    .A(\data_i[16] ),
    .B(_01554_),
    .Y(_04559_)
  );
  AND _12808_ (
    .A(_04558_),
    .B(_04559_),
    .Y(_04560_)
  );
  NAND _12809_ (
    .A(\data_i[8] ),
    .B(_01474_),
    .Y(_04561_)
  );
  AND _12810_ (
    .A(_01470_),
    .B(_04561_),
    .Y(_04562_)
  );
  NAND _12811_ (
    .A(_01475_),
    .B(_04560_),
    .Y(_04563_)
  );
  NAND _12812_ (
    .A(_04562_),
    .B(_04563_),
    .Y(_04564_)
  );
  OR _12813_ (
    .A(\data_i[0] ),
    .B(_01470_),
    .Y(_04565_)
  );
  AND _12814_ (
    .A(MemWrite_i),
    .B(_04565_),
    .Y(_04566_)
  );
  NAND _12815_ (
    .A(_04564_),
    .B(_04566_),
    .Y(_04567_)
  );
  NAND _12816_ (
    .A(_04554_),
    .B(_04567_),
    .Y(_00112_)
  );
  NAND _12817_ (
    .A(\memory[22][1] ),
    .B(_05361_),
    .Y(_04568_)
  );
  OR _12818_ (
    .A(\memory[22][1] ),
    .B(_01534_),
    .Y(_04569_)
  );
  OR _12819_ (
    .A(\data_i[25] ),
    .B(_01535_),
    .Y(_04570_)
  );
  NAND _12820_ (
    .A(_04569_),
    .B(_04570_),
    .Y(_04571_)
  );
  NAND _12821_ (
    .A(_01554_),
    .B(_04571_),
    .Y(_04572_)
  );
  OR _12822_ (
    .A(\data_i[17] ),
    .B(_01554_),
    .Y(_04573_)
  );
  AND _12823_ (
    .A(_04572_),
    .B(_04573_),
    .Y(_04574_)
  );
  NAND _12824_ (
    .A(\data_i[9] ),
    .B(_01474_),
    .Y(_04575_)
  );
  AND _12825_ (
    .A(_01470_),
    .B(_04575_),
    .Y(_04576_)
  );
  NAND _12826_ (
    .A(_01475_),
    .B(_04574_),
    .Y(_04577_)
  );
  NAND _12827_ (
    .A(_04576_),
    .B(_04577_),
    .Y(_04578_)
  );
  OR _12828_ (
    .A(\data_i[1] ),
    .B(_01470_),
    .Y(_04579_)
  );
  AND _12829_ (
    .A(MemWrite_i),
    .B(_04579_),
    .Y(_04580_)
  );
  NAND _12830_ (
    .A(_04578_),
    .B(_04580_),
    .Y(_04581_)
  );
  NAND _12831_ (
    .A(_04568_),
    .B(_04581_),
    .Y(_00113_)
  );
  NAND _12832_ (
    .A(\memory[22][2] ),
    .B(_05361_),
    .Y(_04582_)
  );
  OR _12833_ (
    .A(\memory[22][2] ),
    .B(_01534_),
    .Y(_04583_)
  );
  OR _12834_ (
    .A(\data_i[26] ),
    .B(_01535_),
    .Y(_04584_)
  );
  NAND _12835_ (
    .A(_04583_),
    .B(_04584_),
    .Y(_04585_)
  );
  NAND _12836_ (
    .A(_01554_),
    .B(_04585_),
    .Y(_04586_)
  );
  OR _12837_ (
    .A(\data_i[18] ),
    .B(_01554_),
    .Y(_04587_)
  );
  AND _12838_ (
    .A(_04586_),
    .B(_04587_),
    .Y(_04588_)
  );
  NAND _12839_ (
    .A(\data_i[10] ),
    .B(_01474_),
    .Y(_04589_)
  );
  AND _12840_ (
    .A(_01470_),
    .B(_04589_),
    .Y(_04590_)
  );
  NAND _12841_ (
    .A(_01475_),
    .B(_04588_),
    .Y(_04591_)
  );
  NAND _12842_ (
    .A(_04590_),
    .B(_04591_),
    .Y(_04592_)
  );
  OR _12843_ (
    .A(\data_i[2] ),
    .B(_01470_),
    .Y(_04593_)
  );
  AND _12844_ (
    .A(MemWrite_i),
    .B(_04593_),
    .Y(_04594_)
  );
  NAND _12845_ (
    .A(_04592_),
    .B(_04594_),
    .Y(_04595_)
  );
  NAND _12846_ (
    .A(_04582_),
    .B(_04595_),
    .Y(_00114_)
  );
  NAND _12847_ (
    .A(\memory[22][3] ),
    .B(_05361_),
    .Y(_04596_)
  );
  OR _12848_ (
    .A(\memory[22][3] ),
    .B(_01534_),
    .Y(_04597_)
  );
  OR _12849_ (
    .A(\data_i[27] ),
    .B(_01535_),
    .Y(_04598_)
  );
  NAND _12850_ (
    .A(_04597_),
    .B(_04598_),
    .Y(_04599_)
  );
  NAND _12851_ (
    .A(_01554_),
    .B(_04599_),
    .Y(_04600_)
  );
  OR _12852_ (
    .A(\data_i[19] ),
    .B(_01554_),
    .Y(_04601_)
  );
  AND _12853_ (
    .A(_04600_),
    .B(_04601_),
    .Y(_04602_)
  );
  NAND _12854_ (
    .A(\data_i[11] ),
    .B(_01474_),
    .Y(_04603_)
  );
  AND _12855_ (
    .A(_01470_),
    .B(_04603_),
    .Y(_04604_)
  );
  NAND _12856_ (
    .A(_01475_),
    .B(_04602_),
    .Y(_04605_)
  );
  NAND _12857_ (
    .A(_04604_),
    .B(_04605_),
    .Y(_04606_)
  );
  OR _12858_ (
    .A(\data_i[3] ),
    .B(_01470_),
    .Y(_04607_)
  );
  AND _12859_ (
    .A(MemWrite_i),
    .B(_04607_),
    .Y(_04608_)
  );
  NAND _12860_ (
    .A(_04606_),
    .B(_04608_),
    .Y(_04609_)
  );
  NAND _12861_ (
    .A(_04596_),
    .B(_04609_),
    .Y(_00115_)
  );
  NAND _12862_ (
    .A(\memory[22][4] ),
    .B(_05361_),
    .Y(_04610_)
  );
  OR _12863_ (
    .A(\memory[22][4] ),
    .B(_01534_),
    .Y(_04611_)
  );
  OR _12864_ (
    .A(\data_i[28] ),
    .B(_01535_),
    .Y(_04612_)
  );
  NAND _12865_ (
    .A(_04611_),
    .B(_04612_),
    .Y(_04613_)
  );
  NAND _12866_ (
    .A(_01554_),
    .B(_04613_),
    .Y(_04614_)
  );
  OR _12867_ (
    .A(\data_i[20] ),
    .B(_01554_),
    .Y(_04615_)
  );
  AND _12868_ (
    .A(_04614_),
    .B(_04615_),
    .Y(_04616_)
  );
  NAND _12869_ (
    .A(\data_i[12] ),
    .B(_01474_),
    .Y(_04617_)
  );
  AND _12870_ (
    .A(_01470_),
    .B(_04617_),
    .Y(_04618_)
  );
  NAND _12871_ (
    .A(_01475_),
    .B(_04616_),
    .Y(_04619_)
  );
  NAND _12872_ (
    .A(_04618_),
    .B(_04619_),
    .Y(_04620_)
  );
  OR _12873_ (
    .A(\data_i[4] ),
    .B(_01470_),
    .Y(_04621_)
  );
  AND _12874_ (
    .A(MemWrite_i),
    .B(_04621_),
    .Y(_04622_)
  );
  NAND _12875_ (
    .A(_04620_),
    .B(_04622_),
    .Y(_04623_)
  );
  NAND _12876_ (
    .A(_04610_),
    .B(_04623_),
    .Y(_00116_)
  );
  NAND _12877_ (
    .A(\memory[22][5] ),
    .B(_05361_),
    .Y(_04624_)
  );
  OR _12878_ (
    .A(\memory[22][5] ),
    .B(_01534_),
    .Y(_04625_)
  );
  OR _12879_ (
    .A(\data_i[29] ),
    .B(_01535_),
    .Y(_04626_)
  );
  NAND _12880_ (
    .A(_04625_),
    .B(_04626_),
    .Y(_04627_)
  );
  NAND _12881_ (
    .A(_01554_),
    .B(_04627_),
    .Y(_04628_)
  );
  OR _12882_ (
    .A(\data_i[21] ),
    .B(_01554_),
    .Y(_04629_)
  );
  AND _12883_ (
    .A(_04628_),
    .B(_04629_),
    .Y(_04630_)
  );
  NAND _12884_ (
    .A(\data_i[13] ),
    .B(_01474_),
    .Y(_04631_)
  );
  AND _12885_ (
    .A(_01470_),
    .B(_04631_),
    .Y(_04632_)
  );
  NAND _12886_ (
    .A(_01475_),
    .B(_04630_),
    .Y(_04633_)
  );
  NAND _12887_ (
    .A(_04632_),
    .B(_04633_),
    .Y(_04634_)
  );
  OR _12888_ (
    .A(\data_i[5] ),
    .B(_01470_),
    .Y(_04635_)
  );
  AND _12889_ (
    .A(MemWrite_i),
    .B(_04635_),
    .Y(_04636_)
  );
  NAND _12890_ (
    .A(_04634_),
    .B(_04636_),
    .Y(_04637_)
  );
  NAND _12891_ (
    .A(_04624_),
    .B(_04637_),
    .Y(_00117_)
  );
  NAND _12892_ (
    .A(\memory[22][6] ),
    .B(_05361_),
    .Y(_04638_)
  );
  OR _12893_ (
    .A(\memory[22][6] ),
    .B(_01534_),
    .Y(_04639_)
  );
  OR _12894_ (
    .A(\data_i[30] ),
    .B(_01535_),
    .Y(_04640_)
  );
  NAND _12895_ (
    .A(_04639_),
    .B(_04640_),
    .Y(_04641_)
  );
  NAND _12896_ (
    .A(_01554_),
    .B(_04641_),
    .Y(_04642_)
  );
  OR _12897_ (
    .A(\data_i[22] ),
    .B(_01554_),
    .Y(_04643_)
  );
  AND _12898_ (
    .A(_04642_),
    .B(_04643_),
    .Y(_04644_)
  );
  NAND _12899_ (
    .A(\data_i[14] ),
    .B(_01474_),
    .Y(_04645_)
  );
  AND _12900_ (
    .A(_01470_),
    .B(_04645_),
    .Y(_04646_)
  );
  NAND _12901_ (
    .A(_01475_),
    .B(_04644_),
    .Y(_04647_)
  );
  NAND _12902_ (
    .A(_04646_),
    .B(_04647_),
    .Y(_04648_)
  );
  OR _12903_ (
    .A(\data_i[6] ),
    .B(_01470_),
    .Y(_04649_)
  );
  AND _12904_ (
    .A(MemWrite_i),
    .B(_04649_),
    .Y(_04650_)
  );
  NAND _12905_ (
    .A(_04648_),
    .B(_04650_),
    .Y(_04651_)
  );
  NAND _12906_ (
    .A(_04638_),
    .B(_04651_),
    .Y(_00118_)
  );
  NAND _12907_ (
    .A(\memory[22][7] ),
    .B(_05361_),
    .Y(_04652_)
  );
  OR _12908_ (
    .A(\memory[22][7] ),
    .B(_01534_),
    .Y(_04653_)
  );
  OR _12909_ (
    .A(\data_i[31] ),
    .B(_01535_),
    .Y(_04654_)
  );
  NAND _12910_ (
    .A(_04653_),
    .B(_04654_),
    .Y(_04655_)
  );
  NAND _12911_ (
    .A(_01554_),
    .B(_04655_),
    .Y(_04656_)
  );
  OR _12912_ (
    .A(\data_i[23] ),
    .B(_01554_),
    .Y(_04657_)
  );
  AND _12913_ (
    .A(_04656_),
    .B(_04657_),
    .Y(_04658_)
  );
  NAND _12914_ (
    .A(\data_i[15] ),
    .B(_01474_),
    .Y(_04659_)
  );
  AND _12915_ (
    .A(_01470_),
    .B(_04659_),
    .Y(_04660_)
  );
  NAND _12916_ (
    .A(_01475_),
    .B(_04658_),
    .Y(_04661_)
  );
  NAND _12917_ (
    .A(_04660_),
    .B(_04661_),
    .Y(_04662_)
  );
  OR _12918_ (
    .A(\data_i[7] ),
    .B(_01470_),
    .Y(_04663_)
  );
  AND _12919_ (
    .A(MemWrite_i),
    .B(_04663_),
    .Y(_04664_)
  );
  NAND _12920_ (
    .A(_04662_),
    .B(_04664_),
    .Y(_04665_)
  );
  NAND _12921_ (
    .A(_04652_),
    .B(_04665_),
    .Y(_00119_)
  );
  NAND _12922_ (
    .A(\memory[21][0] ),
    .B(_05361_),
    .Y(_04666_)
  );
  OR _12923_ (
    .A(\memory[21][0] ),
    .B(_01582_),
    .Y(_04667_)
  );
  OR _12924_ (
    .A(\data_i[24] ),
    .B(_01583_),
    .Y(_04668_)
  );
  NAND _12925_ (
    .A(_04667_),
    .B(_04668_),
    .Y(_04669_)
  );
  NAND _12926_ (
    .A(_01535_),
    .B(_04669_),
    .Y(_04670_)
  );
  OR _12927_ (
    .A(\data_i[16] ),
    .B(_01535_),
    .Y(_04671_)
  );
  AND _12928_ (
    .A(_04670_),
    .B(_04671_),
    .Y(_04672_)
  );
  NAND _12929_ (
    .A(\data_i[8] ),
    .B(_01553_),
    .Y(_04673_)
  );
  AND _12930_ (
    .A(_01475_),
    .B(_04673_),
    .Y(_04674_)
  );
  NAND _12931_ (
    .A(_01554_),
    .B(_04672_),
    .Y(_04675_)
  );
  NAND _12932_ (
    .A(_04674_),
    .B(_04675_),
    .Y(_04676_)
  );
  OR _12933_ (
    .A(\data_i[0] ),
    .B(_01475_),
    .Y(_04677_)
  );
  AND _12934_ (
    .A(MemWrite_i),
    .B(_04677_),
    .Y(_04678_)
  );
  NAND _12935_ (
    .A(_04676_),
    .B(_04678_),
    .Y(_04679_)
  );
  NAND _12936_ (
    .A(_04666_),
    .B(_04679_),
    .Y(_00104_)
  );
  NAND _12937_ (
    .A(\memory[21][1] ),
    .B(_05361_),
    .Y(_04680_)
  );
  OR _12938_ (
    .A(\memory[21][1] ),
    .B(_01582_),
    .Y(_04681_)
  );
  OR _12939_ (
    .A(\data_i[25] ),
    .B(_01583_),
    .Y(_04682_)
  );
  NAND _12940_ (
    .A(_04681_),
    .B(_04682_),
    .Y(_04683_)
  );
  NAND _12941_ (
    .A(_01535_),
    .B(_04683_),
    .Y(_04684_)
  );
  OR _12942_ (
    .A(\data_i[17] ),
    .B(_01535_),
    .Y(_04685_)
  );
  AND _12943_ (
    .A(_04684_),
    .B(_04685_),
    .Y(_04686_)
  );
  NAND _12944_ (
    .A(\data_i[9] ),
    .B(_01553_),
    .Y(_04687_)
  );
  AND _12945_ (
    .A(_01475_),
    .B(_04687_),
    .Y(_04688_)
  );
  NAND _12946_ (
    .A(_01554_),
    .B(_04686_),
    .Y(_04689_)
  );
  NAND _12947_ (
    .A(_04688_),
    .B(_04689_),
    .Y(_04690_)
  );
  OR _12948_ (
    .A(\data_i[1] ),
    .B(_01475_),
    .Y(_04691_)
  );
  AND _12949_ (
    .A(MemWrite_i),
    .B(_04691_),
    .Y(_04692_)
  );
  NAND _12950_ (
    .A(_04690_),
    .B(_04692_),
    .Y(_04693_)
  );
  NAND _12951_ (
    .A(_04680_),
    .B(_04693_),
    .Y(_00105_)
  );
  NAND _12952_ (
    .A(\memory[21][2] ),
    .B(_05361_),
    .Y(_04694_)
  );
  OR _12953_ (
    .A(\memory[21][2] ),
    .B(_01582_),
    .Y(_04695_)
  );
  OR _12954_ (
    .A(\data_i[26] ),
    .B(_01583_),
    .Y(_04696_)
  );
  NAND _12955_ (
    .A(_04695_),
    .B(_04696_),
    .Y(_04697_)
  );
  NAND _12956_ (
    .A(_01535_),
    .B(_04697_),
    .Y(_04698_)
  );
  OR _12957_ (
    .A(\data_i[18] ),
    .B(_01535_),
    .Y(_04699_)
  );
  AND _12958_ (
    .A(_04698_),
    .B(_04699_),
    .Y(_04700_)
  );
  NAND _12959_ (
    .A(\data_i[10] ),
    .B(_01553_),
    .Y(_04701_)
  );
  AND _12960_ (
    .A(_01475_),
    .B(_04701_),
    .Y(_04702_)
  );
  NAND _12961_ (
    .A(_01554_),
    .B(_04700_),
    .Y(_04703_)
  );
  NAND _12962_ (
    .A(_04702_),
    .B(_04703_),
    .Y(_04704_)
  );
  OR _12963_ (
    .A(\data_i[2] ),
    .B(_01475_),
    .Y(_04705_)
  );
  AND _12964_ (
    .A(MemWrite_i),
    .B(_04705_),
    .Y(_04706_)
  );
  NAND _12965_ (
    .A(_04704_),
    .B(_04706_),
    .Y(_04707_)
  );
  NAND _12966_ (
    .A(_04694_),
    .B(_04707_),
    .Y(_00106_)
  );
  NAND _12967_ (
    .A(\memory[21][3] ),
    .B(_05361_),
    .Y(_04708_)
  );
  OR _12968_ (
    .A(\memory[21][3] ),
    .B(_01582_),
    .Y(_04709_)
  );
  OR _12969_ (
    .A(\data_i[27] ),
    .B(_01583_),
    .Y(_04710_)
  );
  NAND _12970_ (
    .A(_04709_),
    .B(_04710_),
    .Y(_04711_)
  );
  NAND _12971_ (
    .A(_01535_),
    .B(_04711_),
    .Y(_04712_)
  );
  OR _12972_ (
    .A(\data_i[19] ),
    .B(_01535_),
    .Y(_04713_)
  );
  AND _12973_ (
    .A(_04712_),
    .B(_04713_),
    .Y(_04714_)
  );
  NAND _12974_ (
    .A(\data_i[11] ),
    .B(_01553_),
    .Y(_04715_)
  );
  AND _12975_ (
    .A(_01475_),
    .B(_04715_),
    .Y(_04716_)
  );
  NAND _12976_ (
    .A(_01554_),
    .B(_04714_),
    .Y(_04717_)
  );
  NAND _12977_ (
    .A(_04716_),
    .B(_04717_),
    .Y(_04718_)
  );
  OR _12978_ (
    .A(\data_i[3] ),
    .B(_01475_),
    .Y(_04719_)
  );
  AND _12979_ (
    .A(MemWrite_i),
    .B(_04719_),
    .Y(_04720_)
  );
  NAND _12980_ (
    .A(_04718_),
    .B(_04720_),
    .Y(_04721_)
  );
  NAND _12981_ (
    .A(_04708_),
    .B(_04721_),
    .Y(_00107_)
  );
  NAND _12982_ (
    .A(\memory[21][4] ),
    .B(_05361_),
    .Y(_04722_)
  );
  OR _12983_ (
    .A(\memory[21][4] ),
    .B(_01582_),
    .Y(_04723_)
  );
  OR _12984_ (
    .A(\data_i[28] ),
    .B(_01583_),
    .Y(_04724_)
  );
  NAND _12985_ (
    .A(_04723_),
    .B(_04724_),
    .Y(_04725_)
  );
  NAND _12986_ (
    .A(_01535_),
    .B(_04725_),
    .Y(_04726_)
  );
  OR _12987_ (
    .A(\data_i[20] ),
    .B(_01535_),
    .Y(_04727_)
  );
  AND _12988_ (
    .A(_04726_),
    .B(_04727_),
    .Y(_04728_)
  );
  NAND _12989_ (
    .A(\data_i[12] ),
    .B(_01553_),
    .Y(_04729_)
  );
  AND _12990_ (
    .A(_01475_),
    .B(_04729_),
    .Y(_04730_)
  );
  NAND _12991_ (
    .A(_01554_),
    .B(_04728_),
    .Y(_04731_)
  );
  NAND _12992_ (
    .A(_04730_),
    .B(_04731_),
    .Y(_04732_)
  );
  OR _12993_ (
    .A(\data_i[4] ),
    .B(_01475_),
    .Y(_04733_)
  );
  AND _12994_ (
    .A(MemWrite_i),
    .B(_04733_),
    .Y(_04734_)
  );
  NAND _12995_ (
    .A(_04732_),
    .B(_04734_),
    .Y(_04735_)
  );
  NAND _12996_ (
    .A(_04722_),
    .B(_04735_),
    .Y(_00108_)
  );
  NAND _12997_ (
    .A(\memory[21][5] ),
    .B(_05361_),
    .Y(_04736_)
  );
  OR _12998_ (
    .A(\memory[21][5] ),
    .B(_01582_),
    .Y(_04737_)
  );
  OR _12999_ (
    .A(\data_i[29] ),
    .B(_01583_),
    .Y(_04738_)
  );
  NAND _13000_ (
    .A(_04737_),
    .B(_04738_),
    .Y(_04739_)
  );
  NAND _13001_ (
    .A(_01535_),
    .B(_04739_),
    .Y(_04740_)
  );
  OR _13002_ (
    .A(\data_i[21] ),
    .B(_01535_),
    .Y(_04741_)
  );
  AND _13003_ (
    .A(_04740_),
    .B(_04741_),
    .Y(_04742_)
  );
  NAND _13004_ (
    .A(\data_i[13] ),
    .B(_01553_),
    .Y(_04743_)
  );
  AND _13005_ (
    .A(_01475_),
    .B(_04743_),
    .Y(_04744_)
  );
  NAND _13006_ (
    .A(_01554_),
    .B(_04742_),
    .Y(_04745_)
  );
  NAND _13007_ (
    .A(_04744_),
    .B(_04745_),
    .Y(_04746_)
  );
  OR _13008_ (
    .A(\data_i[5] ),
    .B(_01475_),
    .Y(_04747_)
  );
  AND _13009_ (
    .A(MemWrite_i),
    .B(_04747_),
    .Y(_04748_)
  );
  NAND _13010_ (
    .A(_04746_),
    .B(_04748_),
    .Y(_04749_)
  );
  NAND _13011_ (
    .A(_04736_),
    .B(_04749_),
    .Y(_00109_)
  );
  NAND _13012_ (
    .A(\memory[21][6] ),
    .B(_05361_),
    .Y(_04750_)
  );
  OR _13013_ (
    .A(\memory[21][6] ),
    .B(_01582_),
    .Y(_04751_)
  );
  OR _13014_ (
    .A(\data_i[30] ),
    .B(_01583_),
    .Y(_04752_)
  );
  NAND _13015_ (
    .A(_04751_),
    .B(_04752_),
    .Y(_04753_)
  );
  NAND _13016_ (
    .A(_01535_),
    .B(_04753_),
    .Y(_04754_)
  );
  OR _13017_ (
    .A(\data_i[22] ),
    .B(_01535_),
    .Y(_04755_)
  );
  AND _13018_ (
    .A(_04754_),
    .B(_04755_),
    .Y(_04756_)
  );
  NAND _13019_ (
    .A(\data_i[14] ),
    .B(_01553_),
    .Y(_04757_)
  );
  AND _13020_ (
    .A(_01475_),
    .B(_04757_),
    .Y(_04758_)
  );
  NAND _13021_ (
    .A(_01554_),
    .B(_04756_),
    .Y(_04759_)
  );
  NAND _13022_ (
    .A(_04758_),
    .B(_04759_),
    .Y(_04760_)
  );
  OR _13023_ (
    .A(\data_i[6] ),
    .B(_01475_),
    .Y(_04761_)
  );
  AND _13024_ (
    .A(MemWrite_i),
    .B(_04761_),
    .Y(_04762_)
  );
  NAND _13025_ (
    .A(_04760_),
    .B(_04762_),
    .Y(_04763_)
  );
  NAND _13026_ (
    .A(_04750_),
    .B(_04763_),
    .Y(_00110_)
  );
  NAND _13027_ (
    .A(\memory[21][7] ),
    .B(_05361_),
    .Y(_04764_)
  );
  OR _13028_ (
    .A(\memory[21][7] ),
    .B(_01582_),
    .Y(_04765_)
  );
  OR _13029_ (
    .A(\data_i[31] ),
    .B(_01583_),
    .Y(_04766_)
  );
  NAND _13030_ (
    .A(_04765_),
    .B(_04766_),
    .Y(_04767_)
  );
  NAND _13031_ (
    .A(_01535_),
    .B(_04767_),
    .Y(_04768_)
  );
  OR _13032_ (
    .A(\data_i[23] ),
    .B(_01535_),
    .Y(_04769_)
  );
  AND _13033_ (
    .A(_04768_),
    .B(_04769_),
    .Y(_04770_)
  );
  NAND _13034_ (
    .A(\data_i[15] ),
    .B(_01553_),
    .Y(_04771_)
  );
  AND _13035_ (
    .A(_01475_),
    .B(_04771_),
    .Y(_04772_)
  );
  NAND _13036_ (
    .A(_01554_),
    .B(_04770_),
    .Y(_04773_)
  );
  NAND _13037_ (
    .A(_04772_),
    .B(_04773_),
    .Y(_04774_)
  );
  OR _13038_ (
    .A(\data_i[7] ),
    .B(_01475_),
    .Y(_04775_)
  );
  AND _13039_ (
    .A(MemWrite_i),
    .B(_04775_),
    .Y(_04776_)
  );
  NAND _13040_ (
    .A(_04774_),
    .B(_04776_),
    .Y(_04777_)
  );
  NAND _13041_ (
    .A(_04764_),
    .B(_04777_),
    .Y(_00111_)
  );
  NAND _13042_ (
    .A(\memory[20][0] ),
    .B(_05361_),
    .Y(_04778_)
  );
  OR _13043_ (
    .A(\memory[20][0] ),
    .B(_01479_),
    .Y(_04779_)
  );
  OR _13044_ (
    .A(\data_i[24] ),
    .B(_01480_),
    .Y(_04780_)
  );
  NAND _13045_ (
    .A(_04779_),
    .B(_04780_),
    .Y(_04781_)
  );
  NAND _13046_ (
    .A(_01583_),
    .B(_04781_),
    .Y(_04782_)
  );
  OR _13047_ (
    .A(\data_i[16] ),
    .B(_01583_),
    .Y(_04783_)
  );
  AND _13048_ (
    .A(_04782_),
    .B(_04783_),
    .Y(_04784_)
  );
  NAND _13049_ (
    .A(\data_i[8] ),
    .B(_01534_),
    .Y(_04785_)
  );
  AND _13050_ (
    .A(_01554_),
    .B(_04785_),
    .Y(_04786_)
  );
  NAND _13051_ (
    .A(_01535_),
    .B(_04784_),
    .Y(_04787_)
  );
  NAND _13052_ (
    .A(_04786_),
    .B(_04787_),
    .Y(_04788_)
  );
  OR _13053_ (
    .A(\data_i[0] ),
    .B(_01554_),
    .Y(_04789_)
  );
  AND _13054_ (
    .A(MemWrite_i),
    .B(_04789_),
    .Y(_04790_)
  );
  NAND _13055_ (
    .A(_04788_),
    .B(_04790_),
    .Y(_04791_)
  );
  NAND _13056_ (
    .A(_04778_),
    .B(_04791_),
    .Y(_00096_)
  );
  NAND _13057_ (
    .A(\memory[20][1] ),
    .B(_05361_),
    .Y(_04792_)
  );
  OR _13058_ (
    .A(\memory[20][1] ),
    .B(_01479_),
    .Y(_04793_)
  );
  OR _13059_ (
    .A(\data_i[25] ),
    .B(_01480_),
    .Y(_04794_)
  );
  NAND _13060_ (
    .A(_04793_),
    .B(_04794_),
    .Y(_04795_)
  );
  NAND _13061_ (
    .A(_01583_),
    .B(_04795_),
    .Y(_04796_)
  );
  OR _13062_ (
    .A(\data_i[17] ),
    .B(_01583_),
    .Y(_04797_)
  );
  AND _13063_ (
    .A(_04796_),
    .B(_04797_),
    .Y(_04798_)
  );
  NAND _13064_ (
    .A(\data_i[9] ),
    .B(_01534_),
    .Y(_04799_)
  );
  AND _13065_ (
    .A(_01554_),
    .B(_04799_),
    .Y(_04800_)
  );
  NAND _13066_ (
    .A(_01535_),
    .B(_04798_),
    .Y(_04801_)
  );
  NAND _13067_ (
    .A(_04800_),
    .B(_04801_),
    .Y(_04802_)
  );
  OR _13068_ (
    .A(\data_i[1] ),
    .B(_01554_),
    .Y(_04803_)
  );
  AND _13069_ (
    .A(MemWrite_i),
    .B(_04803_),
    .Y(_04804_)
  );
  NAND _13070_ (
    .A(_04802_),
    .B(_04804_),
    .Y(_04805_)
  );
  NAND _13071_ (
    .A(_04792_),
    .B(_04805_),
    .Y(_00097_)
  );
  OR _13072_ (
    .A(\memory[20][2] ),
    .B(MemWrite_i),
    .Y(_04806_)
  );
  NAND _13073_ (
    .A(\data_i[26] ),
    .B(_01479_),
    .Y(_04807_)
  );
  NAND _13074_ (
    .A(\memory[20][2] ),
    .B(_01480_),
    .Y(_04808_)
  );
  NAND _13075_ (
    .A(_04807_),
    .B(_04808_),
    .Y(_04809_)
  );
  NAND _13076_ (
    .A(_01583_),
    .B(_04809_),
    .Y(_04810_)
  );
  NAND _13077_ (
    .A(\data_i[18] ),
    .B(_01582_),
    .Y(_04811_)
  );
  AND _13078_ (
    .A(_01535_),
    .B(_04811_),
    .Y(_04812_)
  );
  NAND _13079_ (
    .A(_04810_),
    .B(_04812_),
    .Y(_04813_)
  );
  OR _13080_ (
    .A(\data_i[10] ),
    .B(_01535_),
    .Y(_04814_)
  );
  AND _13081_ (
    .A(_01554_),
    .B(_04814_),
    .Y(_04815_)
  );
  NAND _13082_ (
    .A(_04813_),
    .B(_04815_),
    .Y(_04816_)
  );
  NAND _13083_ (
    .A(\data_i[2] ),
    .B(_01553_),
    .Y(_04817_)
  );
  AND _13084_ (
    .A(MemWrite_i),
    .B(_04817_),
    .Y(_04818_)
  );
  NAND _13085_ (
    .A(_04816_),
    .B(_04818_),
    .Y(_04819_)
  );
  AND _13086_ (
    .A(_04806_),
    .B(_04819_),
    .Y(_00098_)
  );
  OR _13087_ (
    .A(\memory[20][3] ),
    .B(MemWrite_i),
    .Y(_04820_)
  );
  NAND _13088_ (
    .A(\data_i[27] ),
    .B(_01479_),
    .Y(_04821_)
  );
  NAND _13089_ (
    .A(\memory[20][3] ),
    .B(_01480_),
    .Y(_04822_)
  );
  NAND _13090_ (
    .A(_04821_),
    .B(_04822_),
    .Y(_04823_)
  );
  NAND _13091_ (
    .A(_01583_),
    .B(_04823_),
    .Y(_04824_)
  );
  NAND _13092_ (
    .A(\data_i[19] ),
    .B(_01582_),
    .Y(_04825_)
  );
  AND _13093_ (
    .A(_01535_),
    .B(_04825_),
    .Y(_04826_)
  );
  NAND _13094_ (
    .A(_04824_),
    .B(_04826_),
    .Y(_04827_)
  );
  OR _13095_ (
    .A(\data_i[11] ),
    .B(_01535_),
    .Y(_04828_)
  );
  AND _13096_ (
    .A(_01554_),
    .B(_04828_),
    .Y(_04829_)
  );
  NAND _13097_ (
    .A(_04827_),
    .B(_04829_),
    .Y(_04830_)
  );
  NAND _13098_ (
    .A(\data_i[3] ),
    .B(_01553_),
    .Y(_04831_)
  );
  AND _13099_ (
    .A(MemWrite_i),
    .B(_04831_),
    .Y(_04832_)
  );
  NAND _13100_ (
    .A(_04830_),
    .B(_04832_),
    .Y(_04833_)
  );
  AND _13101_ (
    .A(_04820_),
    .B(_04833_),
    .Y(_00099_)
  );
  OR _13102_ (
    .A(\memory[20][4] ),
    .B(MemWrite_i),
    .Y(_04834_)
  );
  NAND _13103_ (
    .A(\data_i[28] ),
    .B(_01479_),
    .Y(_04835_)
  );
  NAND _13104_ (
    .A(\memory[20][4] ),
    .B(_01480_),
    .Y(_04836_)
  );
  NAND _13105_ (
    .A(_04835_),
    .B(_04836_),
    .Y(_04837_)
  );
  NAND _13106_ (
    .A(_01583_),
    .B(_04837_),
    .Y(_04838_)
  );
  NAND _13107_ (
    .A(\data_i[20] ),
    .B(_01582_),
    .Y(_04839_)
  );
  AND _13108_ (
    .A(_01535_),
    .B(_04839_),
    .Y(_04840_)
  );
  NAND _13109_ (
    .A(_04838_),
    .B(_04840_),
    .Y(_04841_)
  );
  OR _13110_ (
    .A(\data_i[12] ),
    .B(_01535_),
    .Y(_04842_)
  );
  AND _13111_ (
    .A(_01554_),
    .B(_04842_),
    .Y(_04843_)
  );
  NAND _13112_ (
    .A(_04841_),
    .B(_04843_),
    .Y(_04844_)
  );
  NAND _13113_ (
    .A(\data_i[4] ),
    .B(_01553_),
    .Y(_04845_)
  );
  AND _13114_ (
    .A(MemWrite_i),
    .B(_04845_),
    .Y(_04846_)
  );
  NAND _13115_ (
    .A(_04844_),
    .B(_04846_),
    .Y(_04847_)
  );
  AND _13116_ (
    .A(_04834_),
    .B(_04847_),
    .Y(_00100_)
  );
  NAND _13117_ (
    .A(\memory[20][5] ),
    .B(_05361_),
    .Y(_04848_)
  );
  OR _13118_ (
    .A(\memory[20][5] ),
    .B(_01479_),
    .Y(_04849_)
  );
  OR _13119_ (
    .A(\data_i[29] ),
    .B(_01480_),
    .Y(_04850_)
  );
  NAND _13120_ (
    .A(_04849_),
    .B(_04850_),
    .Y(_04851_)
  );
  NAND _13121_ (
    .A(_01583_),
    .B(_04851_),
    .Y(_04852_)
  );
  OR _13122_ (
    .A(\data_i[21] ),
    .B(_01583_),
    .Y(_04853_)
  );
  AND _13123_ (
    .A(_04852_),
    .B(_04853_),
    .Y(_04854_)
  );
  NAND _13124_ (
    .A(\data_i[13] ),
    .B(_01534_),
    .Y(_04855_)
  );
  AND _13125_ (
    .A(_01554_),
    .B(_04855_),
    .Y(_04856_)
  );
  NAND _13126_ (
    .A(_01535_),
    .B(_04854_),
    .Y(_04857_)
  );
  NAND _13127_ (
    .A(_04856_),
    .B(_04857_),
    .Y(_04858_)
  );
  OR _13128_ (
    .A(\data_i[5] ),
    .B(_01554_),
    .Y(_04859_)
  );
  AND _13129_ (
    .A(MemWrite_i),
    .B(_04859_),
    .Y(_04860_)
  );
  NAND _13130_ (
    .A(_04858_),
    .B(_04860_),
    .Y(_04861_)
  );
  NAND _13131_ (
    .A(_04848_),
    .B(_04861_),
    .Y(_00101_)
  );
  NAND _13132_ (
    .A(\memory[20][6] ),
    .B(_05361_),
    .Y(_04862_)
  );
  OR _13133_ (
    .A(\memory[20][6] ),
    .B(_01479_),
    .Y(_04863_)
  );
  OR _13134_ (
    .A(\data_i[30] ),
    .B(_01480_),
    .Y(_04864_)
  );
  NAND _13135_ (
    .A(_04863_),
    .B(_04864_),
    .Y(_04865_)
  );
  NAND _13136_ (
    .A(_01583_),
    .B(_04865_),
    .Y(_04866_)
  );
  OR _13137_ (
    .A(\data_i[22] ),
    .B(_01583_),
    .Y(_04867_)
  );
  AND _13138_ (
    .A(_04866_),
    .B(_04867_),
    .Y(_04868_)
  );
  NAND _13139_ (
    .A(\data_i[14] ),
    .B(_01534_),
    .Y(_04869_)
  );
  AND _13140_ (
    .A(_01554_),
    .B(_04869_),
    .Y(_04870_)
  );
  NAND _13141_ (
    .A(_01535_),
    .B(_04868_),
    .Y(_04871_)
  );
  NAND _13142_ (
    .A(_04870_),
    .B(_04871_),
    .Y(_04872_)
  );
  OR _13143_ (
    .A(\data_i[6] ),
    .B(_01554_),
    .Y(_04873_)
  );
  AND _13144_ (
    .A(MemWrite_i),
    .B(_04873_),
    .Y(_04874_)
  );
  NAND _13145_ (
    .A(_04872_),
    .B(_04874_),
    .Y(_04875_)
  );
  NAND _13146_ (
    .A(_04862_),
    .B(_04875_),
    .Y(_00102_)
  );
  NAND _13147_ (
    .A(\memory[20][7] ),
    .B(_05361_),
    .Y(_04876_)
  );
  OR _13148_ (
    .A(\memory[20][7] ),
    .B(_01479_),
    .Y(_04877_)
  );
  OR _13149_ (
    .A(\data_i[31] ),
    .B(_01480_),
    .Y(_04878_)
  );
  NAND _13150_ (
    .A(_04877_),
    .B(_04878_),
    .Y(_04879_)
  );
  NAND _13151_ (
    .A(_01583_),
    .B(_04879_),
    .Y(_04880_)
  );
  OR _13152_ (
    .A(\data_i[23] ),
    .B(_01583_),
    .Y(_04881_)
  );
  AND _13153_ (
    .A(_04880_),
    .B(_04881_),
    .Y(_04882_)
  );
  NAND _13154_ (
    .A(\data_i[15] ),
    .B(_01534_),
    .Y(_04883_)
  );
  AND _13155_ (
    .A(_01554_),
    .B(_04883_),
    .Y(_04884_)
  );
  NAND _13156_ (
    .A(_01535_),
    .B(_04882_),
    .Y(_04885_)
  );
  NAND _13157_ (
    .A(_04884_),
    .B(_04885_),
    .Y(_04886_)
  );
  OR _13158_ (
    .A(\data_i[7] ),
    .B(_01554_),
    .Y(_04887_)
  );
  AND _13159_ (
    .A(MemWrite_i),
    .B(_04887_),
    .Y(_04888_)
  );
  NAND _13160_ (
    .A(_04886_),
    .B(_04888_),
    .Y(_04889_)
  );
  NAND _13161_ (
    .A(_04876_),
    .B(_04889_),
    .Y(_00103_)
  );
  NAND _13162_ (
    .A(\memory[19][0] ),
    .B(_05361_),
    .Y(_04890_)
  );
  OR _13163_ (
    .A(\memory[19][0] ),
    .B(_01567_),
    .Y(_04891_)
  );
  OR _13164_ (
    .A(\data_i[24] ),
    .B(_01568_),
    .Y(_04892_)
  );
  NAND _13165_ (
    .A(_04891_),
    .B(_04892_),
    .Y(_04893_)
  );
  NAND _13166_ (
    .A(_01480_),
    .B(_04893_),
    .Y(_04894_)
  );
  OR _13167_ (
    .A(\data_i[16] ),
    .B(_01480_),
    .Y(_04895_)
  );
  AND _13168_ (
    .A(_04894_),
    .B(_04895_),
    .Y(_04896_)
  );
  NAND _13169_ (
    .A(\data_i[8] ),
    .B(_01582_),
    .Y(_04897_)
  );
  AND _13170_ (
    .A(_01535_),
    .B(_04897_),
    .Y(_04898_)
  );
  NAND _13171_ (
    .A(_01583_),
    .B(_04896_),
    .Y(_04899_)
  );
  NAND _13172_ (
    .A(_04898_),
    .B(_04899_),
    .Y(_04900_)
  );
  OR _13173_ (
    .A(\data_i[0] ),
    .B(_01535_),
    .Y(_04901_)
  );
  AND _13174_ (
    .A(MemWrite_i),
    .B(_04901_),
    .Y(_04902_)
  );
  NAND _13175_ (
    .A(_04900_),
    .B(_04902_),
    .Y(_04903_)
  );
  NAND _13176_ (
    .A(_04890_),
    .B(_04903_),
    .Y(_00080_)
  );
  NAND _13177_ (
    .A(\memory[19][1] ),
    .B(_05361_),
    .Y(_04904_)
  );
  OR _13178_ (
    .A(\memory[19][1] ),
    .B(_01567_),
    .Y(_04905_)
  );
  OR _13179_ (
    .A(\data_i[25] ),
    .B(_01568_),
    .Y(_04906_)
  );
  NAND _13180_ (
    .A(_04905_),
    .B(_04906_),
    .Y(_04907_)
  );
  NAND _13181_ (
    .A(_01480_),
    .B(_04907_),
    .Y(_04908_)
  );
  OR _13182_ (
    .A(\data_i[17] ),
    .B(_01480_),
    .Y(_04909_)
  );
  AND _13183_ (
    .A(_04908_),
    .B(_04909_),
    .Y(_04910_)
  );
  NAND _13184_ (
    .A(\data_i[9] ),
    .B(_01582_),
    .Y(_04911_)
  );
  AND _13185_ (
    .A(_01535_),
    .B(_04911_),
    .Y(_04912_)
  );
  NAND _13186_ (
    .A(_01583_),
    .B(_04910_),
    .Y(_04913_)
  );
  NAND _13187_ (
    .A(_04912_),
    .B(_04913_),
    .Y(_04914_)
  );
  OR _13188_ (
    .A(\data_i[1] ),
    .B(_01535_),
    .Y(_04915_)
  );
  AND _13189_ (
    .A(MemWrite_i),
    .B(_04915_),
    .Y(_04916_)
  );
  NAND _13190_ (
    .A(_04914_),
    .B(_04916_),
    .Y(_04917_)
  );
  NAND _13191_ (
    .A(_04904_),
    .B(_04917_),
    .Y(_00081_)
  );
  NAND _13192_ (
    .A(\memory[19][2] ),
    .B(_05361_),
    .Y(_04918_)
  );
  OR _13193_ (
    .A(\memory[19][2] ),
    .B(_01567_),
    .Y(_04919_)
  );
  OR _13194_ (
    .A(\data_i[26] ),
    .B(_01568_),
    .Y(_04920_)
  );
  NAND _13195_ (
    .A(_04919_),
    .B(_04920_),
    .Y(_04921_)
  );
  NAND _13196_ (
    .A(_01480_),
    .B(_04921_),
    .Y(_04922_)
  );
  OR _13197_ (
    .A(\data_i[18] ),
    .B(_01480_),
    .Y(_04923_)
  );
  AND _13198_ (
    .A(_04922_),
    .B(_04923_),
    .Y(_04924_)
  );
  NAND _13199_ (
    .A(\data_i[10] ),
    .B(_01582_),
    .Y(_04925_)
  );
  AND _13200_ (
    .A(_01535_),
    .B(_04925_),
    .Y(_04926_)
  );
  NAND _13201_ (
    .A(_01583_),
    .B(_04924_),
    .Y(_04927_)
  );
  NAND _13202_ (
    .A(_04926_),
    .B(_04927_),
    .Y(_04928_)
  );
  OR _13203_ (
    .A(\data_i[2] ),
    .B(_01535_),
    .Y(_04929_)
  );
  AND _13204_ (
    .A(MemWrite_i),
    .B(_04929_),
    .Y(_04930_)
  );
  NAND _13205_ (
    .A(_04928_),
    .B(_04930_),
    .Y(_04931_)
  );
  NAND _13206_ (
    .A(_04918_),
    .B(_04931_),
    .Y(_00082_)
  );
  NAND _13207_ (
    .A(\memory[19][3] ),
    .B(_05361_),
    .Y(_04932_)
  );
  OR _13208_ (
    .A(\memory[19][3] ),
    .B(_01567_),
    .Y(_04933_)
  );
  OR _13209_ (
    .A(\data_i[27] ),
    .B(_01568_),
    .Y(_04934_)
  );
  NAND _13210_ (
    .A(_04933_),
    .B(_04934_),
    .Y(_04935_)
  );
  NAND _13211_ (
    .A(_01480_),
    .B(_04935_),
    .Y(_04936_)
  );
  OR _13212_ (
    .A(\data_i[19] ),
    .B(_01480_),
    .Y(_04937_)
  );
  AND _13213_ (
    .A(_04936_),
    .B(_04937_),
    .Y(_04938_)
  );
  NAND _13214_ (
    .A(\data_i[11] ),
    .B(_01582_),
    .Y(_04939_)
  );
  AND _13215_ (
    .A(_01535_),
    .B(_04939_),
    .Y(_04940_)
  );
  NAND _13216_ (
    .A(_01583_),
    .B(_04938_),
    .Y(_04941_)
  );
  NAND _13217_ (
    .A(_04940_),
    .B(_04941_),
    .Y(_04942_)
  );
  OR _13218_ (
    .A(\data_i[3] ),
    .B(_01535_),
    .Y(_04943_)
  );
  AND _13219_ (
    .A(MemWrite_i),
    .B(_04943_),
    .Y(_04944_)
  );
  NAND _13220_ (
    .A(_04942_),
    .B(_04944_),
    .Y(_04945_)
  );
  NAND _13221_ (
    .A(_04932_),
    .B(_04945_),
    .Y(_00083_)
  );
  OR _13222_ (
    .A(\memory[19][4] ),
    .B(MemWrite_i),
    .Y(_04946_)
  );
  NAND _13223_ (
    .A(\data_i[28] ),
    .B(_01567_),
    .Y(_04947_)
  );
  NAND _13224_ (
    .A(\memory[19][4] ),
    .B(_01568_),
    .Y(_04948_)
  );
  NAND _13225_ (
    .A(_04947_),
    .B(_04948_),
    .Y(_04949_)
  );
  NAND _13226_ (
    .A(_01480_),
    .B(_04949_),
    .Y(_04950_)
  );
  NAND _13227_ (
    .A(\data_i[20] ),
    .B(_01479_),
    .Y(_04951_)
  );
  AND _13228_ (
    .A(_01583_),
    .B(_04951_),
    .Y(_04952_)
  );
  NAND _13229_ (
    .A(_04950_),
    .B(_04952_),
    .Y(_04953_)
  );
  OR _13230_ (
    .A(\data_i[12] ),
    .B(_01583_),
    .Y(_04954_)
  );
  AND _13231_ (
    .A(_01535_),
    .B(_04954_),
    .Y(_04955_)
  );
  NAND _13232_ (
    .A(_04953_),
    .B(_04955_),
    .Y(_04956_)
  );
  NAND _13233_ (
    .A(\data_i[4] ),
    .B(_01534_),
    .Y(_04957_)
  );
  AND _13234_ (
    .A(MemWrite_i),
    .B(_04957_),
    .Y(_04958_)
  );
  NAND _13235_ (
    .A(_04956_),
    .B(_04958_),
    .Y(_04959_)
  );
  AND _13236_ (
    .A(_04946_),
    .B(_04959_),
    .Y(_00084_)
  );
  NAND _13237_ (
    .A(\memory[19][5] ),
    .B(_05361_),
    .Y(_04960_)
  );
  OR _13238_ (
    .A(\memory[19][5] ),
    .B(_01567_),
    .Y(_04961_)
  );
  OR _13239_ (
    .A(\data_i[29] ),
    .B(_01568_),
    .Y(_04962_)
  );
  NAND _13240_ (
    .A(_04961_),
    .B(_04962_),
    .Y(_04963_)
  );
  NAND _13241_ (
    .A(_01480_),
    .B(_04963_),
    .Y(_04964_)
  );
  OR _13242_ (
    .A(\data_i[21] ),
    .B(_01480_),
    .Y(_04965_)
  );
  AND _13243_ (
    .A(_04964_),
    .B(_04965_),
    .Y(_04966_)
  );
  NAND _13244_ (
    .A(\data_i[13] ),
    .B(_01582_),
    .Y(_04967_)
  );
  AND _13245_ (
    .A(_01535_),
    .B(_04967_),
    .Y(_04968_)
  );
  NAND _13246_ (
    .A(_01583_),
    .B(_04966_),
    .Y(_04969_)
  );
  NAND _13247_ (
    .A(_04968_),
    .B(_04969_),
    .Y(_04970_)
  );
  OR _13248_ (
    .A(\data_i[5] ),
    .B(_01535_),
    .Y(_04971_)
  );
  AND _13249_ (
    .A(MemWrite_i),
    .B(_04971_),
    .Y(_04972_)
  );
  NAND _13250_ (
    .A(_04970_),
    .B(_04972_),
    .Y(_04973_)
  );
  NAND _13251_ (
    .A(_04960_),
    .B(_04973_),
    .Y(_00085_)
  );
  OR _13252_ (
    .A(\memory[19][6] ),
    .B(MemWrite_i),
    .Y(_04974_)
  );
  NAND _13253_ (
    .A(\data_i[30] ),
    .B(_01567_),
    .Y(_04975_)
  );
  NAND _13254_ (
    .A(\memory[19][6] ),
    .B(_01568_),
    .Y(_04976_)
  );
  NAND _13255_ (
    .A(_04975_),
    .B(_04976_),
    .Y(_04977_)
  );
  NAND _13256_ (
    .A(_01480_),
    .B(_04977_),
    .Y(_04978_)
  );
  NAND _13257_ (
    .A(\data_i[22] ),
    .B(_01479_),
    .Y(_04979_)
  );
  AND _13258_ (
    .A(_01583_),
    .B(_04979_),
    .Y(_04980_)
  );
  NAND _13259_ (
    .A(_04978_),
    .B(_04980_),
    .Y(_04981_)
  );
  OR _13260_ (
    .A(\data_i[14] ),
    .B(_01583_),
    .Y(_04982_)
  );
  AND _13261_ (
    .A(_01535_),
    .B(_04982_),
    .Y(_04983_)
  );
  NAND _13262_ (
    .A(_04981_),
    .B(_04983_),
    .Y(_04984_)
  );
  NAND _13263_ (
    .A(\data_i[6] ),
    .B(_01534_),
    .Y(_04985_)
  );
  AND _13264_ (
    .A(MemWrite_i),
    .B(_04985_),
    .Y(_04986_)
  );
  NAND _13265_ (
    .A(_04984_),
    .B(_04986_),
    .Y(_04987_)
  );
  AND _13266_ (
    .A(_04974_),
    .B(_04987_),
    .Y(_00086_)
  );
  NAND _13267_ (
    .A(\memory[19][7] ),
    .B(_05361_),
    .Y(_04988_)
  );
  OR _13268_ (
    .A(\memory[19][7] ),
    .B(_01567_),
    .Y(_04989_)
  );
  OR _13269_ (
    .A(\data_i[31] ),
    .B(_01568_),
    .Y(_04990_)
  );
  NAND _13270_ (
    .A(_04989_),
    .B(_04990_),
    .Y(_04991_)
  );
  NAND _13271_ (
    .A(_01480_),
    .B(_04991_),
    .Y(_04992_)
  );
  OR _13272_ (
    .A(\data_i[23] ),
    .B(_01480_),
    .Y(_04993_)
  );
  AND _13273_ (
    .A(_04992_),
    .B(_04993_),
    .Y(_04994_)
  );
  NAND _13274_ (
    .A(\data_i[15] ),
    .B(_01582_),
    .Y(_04995_)
  );
  AND _13275_ (
    .A(_01535_),
    .B(_04995_),
    .Y(_04996_)
  );
  NAND _13276_ (
    .A(_01583_),
    .B(_04994_),
    .Y(_04997_)
  );
  NAND _13277_ (
    .A(_04996_),
    .B(_04997_),
    .Y(_04998_)
  );
  OR _13278_ (
    .A(\data_i[7] ),
    .B(_01535_),
    .Y(_04999_)
  );
  AND _13279_ (
    .A(MemWrite_i),
    .B(_04999_),
    .Y(_05000_)
  );
  NAND _13280_ (
    .A(_04998_),
    .B(_05000_),
    .Y(_05001_)
  );
  NAND _13281_ (
    .A(_04988_),
    .B(_05001_),
    .Y(_00087_)
  );
  NAND _13282_ (
    .A(\memory[18][0] ),
    .B(_05361_),
    .Y(_05002_)
  );
  OR _13283_ (
    .A(\memory[18][0] ),
    .B(_01501_),
    .Y(_05003_)
  );
  OR _13284_ (
    .A(\data_i[24] ),
    .B(_01502_),
    .Y(_05004_)
  );
  NAND _13285_ (
    .A(_05003_),
    .B(_05004_),
    .Y(_05005_)
  );
  NAND _13286_ (
    .A(_01568_),
    .B(_05005_),
    .Y(_05006_)
  );
  OR _13287_ (
    .A(\data_i[16] ),
    .B(_01568_),
    .Y(_05007_)
  );
  AND _13288_ (
    .A(_05006_),
    .B(_05007_),
    .Y(_05008_)
  );
  NAND _13289_ (
    .A(\data_i[8] ),
    .B(_01479_),
    .Y(_05009_)
  );
  AND _13290_ (
    .A(_01583_),
    .B(_05009_),
    .Y(_05010_)
  );
  NAND _13291_ (
    .A(_01480_),
    .B(_05008_),
    .Y(_05011_)
  );
  NAND _13292_ (
    .A(_05010_),
    .B(_05011_),
    .Y(_05012_)
  );
  OR _13293_ (
    .A(\data_i[0] ),
    .B(_01583_),
    .Y(_05013_)
  );
  AND _13294_ (
    .A(MemWrite_i),
    .B(_05013_),
    .Y(_05014_)
  );
  NAND _13295_ (
    .A(_05012_),
    .B(_05014_),
    .Y(_05015_)
  );
  NAND _13296_ (
    .A(_05002_),
    .B(_05015_),
    .Y(_00072_)
  );
  NAND _13297_ (
    .A(\memory[18][1] ),
    .B(_05361_),
    .Y(_05016_)
  );
  OR _13298_ (
    .A(\memory[18][1] ),
    .B(_01501_),
    .Y(_05017_)
  );
  OR _13299_ (
    .A(\data_i[25] ),
    .B(_01502_),
    .Y(_05018_)
  );
  NAND _13300_ (
    .A(_05017_),
    .B(_05018_),
    .Y(_05019_)
  );
  NAND _13301_ (
    .A(_01568_),
    .B(_05019_),
    .Y(_05020_)
  );
  OR _13302_ (
    .A(\data_i[17] ),
    .B(_01568_),
    .Y(_05021_)
  );
  AND _13303_ (
    .A(_05020_),
    .B(_05021_),
    .Y(_05022_)
  );
  NAND _13304_ (
    .A(\data_i[9] ),
    .B(_01479_),
    .Y(_05023_)
  );
  AND _13305_ (
    .A(_01583_),
    .B(_05023_),
    .Y(_05024_)
  );
  NAND _13306_ (
    .A(_01480_),
    .B(_05022_),
    .Y(_05025_)
  );
  NAND _13307_ (
    .A(_05024_),
    .B(_05025_),
    .Y(_05026_)
  );
  OR _13308_ (
    .A(\data_i[1] ),
    .B(_01583_),
    .Y(_05027_)
  );
  AND _13309_ (
    .A(MemWrite_i),
    .B(_05027_),
    .Y(_05028_)
  );
  NAND _13310_ (
    .A(_05026_),
    .B(_05028_),
    .Y(_05029_)
  );
  NAND _13311_ (
    .A(_05016_),
    .B(_05029_),
    .Y(_00073_)
  );
  NAND _13312_ (
    .A(\memory[18][2] ),
    .B(_05361_),
    .Y(_05030_)
  );
  OR _13313_ (
    .A(\memory[18][2] ),
    .B(_01501_),
    .Y(_05031_)
  );
  OR _13314_ (
    .A(\data_i[26] ),
    .B(_01502_),
    .Y(_05032_)
  );
  NAND _13315_ (
    .A(_05031_),
    .B(_05032_),
    .Y(_05033_)
  );
  NAND _13316_ (
    .A(_01568_),
    .B(_05033_),
    .Y(_05034_)
  );
  OR _13317_ (
    .A(\data_i[18] ),
    .B(_01568_),
    .Y(_05035_)
  );
  AND _13318_ (
    .A(_05034_),
    .B(_05035_),
    .Y(_05036_)
  );
  NAND _13319_ (
    .A(\data_i[10] ),
    .B(_01479_),
    .Y(_05037_)
  );
  AND _13320_ (
    .A(_01583_),
    .B(_05037_),
    .Y(_05038_)
  );
  NAND _13321_ (
    .A(_01480_),
    .B(_05036_),
    .Y(_05039_)
  );
  NAND _13322_ (
    .A(_05038_),
    .B(_05039_),
    .Y(_05040_)
  );
  OR _13323_ (
    .A(\data_i[2] ),
    .B(_01583_),
    .Y(_05041_)
  );
  AND _13324_ (
    .A(MemWrite_i),
    .B(_05041_),
    .Y(_05042_)
  );
  NAND _13325_ (
    .A(_05040_),
    .B(_05042_),
    .Y(_05043_)
  );
  NAND _13326_ (
    .A(_05030_),
    .B(_05043_),
    .Y(_00074_)
  );
  OR _13327_ (
    .A(\memory[18][3] ),
    .B(MemWrite_i),
    .Y(_05044_)
  );
  NAND _13328_ (
    .A(\data_i[27] ),
    .B(_01501_),
    .Y(_05045_)
  );
  NAND _13329_ (
    .A(\memory[18][3] ),
    .B(_01502_),
    .Y(_05046_)
  );
  NAND _13330_ (
    .A(_05045_),
    .B(_05046_),
    .Y(_05047_)
  );
  NAND _13331_ (
    .A(_01568_),
    .B(_05047_),
    .Y(_05048_)
  );
  NAND _13332_ (
    .A(\data_i[19] ),
    .B(_01567_),
    .Y(_05049_)
  );
  AND _13333_ (
    .A(_01480_),
    .B(_05049_),
    .Y(_05050_)
  );
  NAND _13334_ (
    .A(_05048_),
    .B(_05050_),
    .Y(_05051_)
  );
  OR _13335_ (
    .A(\data_i[11] ),
    .B(_01480_),
    .Y(_05052_)
  );
  AND _13336_ (
    .A(_01583_),
    .B(_05052_),
    .Y(_05053_)
  );
  NAND _13337_ (
    .A(_05051_),
    .B(_05053_),
    .Y(_05054_)
  );
  NAND _13338_ (
    .A(\data_i[3] ),
    .B(_01582_),
    .Y(_05055_)
  );
  AND _13339_ (
    .A(MemWrite_i),
    .B(_05055_),
    .Y(_05056_)
  );
  NAND _13340_ (
    .A(_05054_),
    .B(_05056_),
    .Y(_05057_)
  );
  AND _13341_ (
    .A(_05044_),
    .B(_05057_),
    .Y(_00075_)
  );
  NAND _13342_ (
    .A(\memory[18][4] ),
    .B(_05361_),
    .Y(_05058_)
  );
  OR _13343_ (
    .A(\memory[18][4] ),
    .B(_01501_),
    .Y(_05059_)
  );
  OR _13344_ (
    .A(\data_i[28] ),
    .B(_01502_),
    .Y(_05060_)
  );
  NAND _13345_ (
    .A(_05059_),
    .B(_05060_),
    .Y(_05061_)
  );
  NAND _13346_ (
    .A(_01568_),
    .B(_05061_),
    .Y(_05062_)
  );
  OR _13347_ (
    .A(\data_i[20] ),
    .B(_01568_),
    .Y(_05063_)
  );
  AND _13348_ (
    .A(_05062_),
    .B(_05063_),
    .Y(_05064_)
  );
  NAND _13349_ (
    .A(\data_i[12] ),
    .B(_01479_),
    .Y(_05065_)
  );
  AND _13350_ (
    .A(_01583_),
    .B(_05065_),
    .Y(_05066_)
  );
  NAND _13351_ (
    .A(_01480_),
    .B(_05064_),
    .Y(_05067_)
  );
  NAND _13352_ (
    .A(_05066_),
    .B(_05067_),
    .Y(_05068_)
  );
  OR _13353_ (
    .A(\data_i[4] ),
    .B(_01583_),
    .Y(_05069_)
  );
  AND _13354_ (
    .A(MemWrite_i),
    .B(_05069_),
    .Y(_05070_)
  );
  NAND _13355_ (
    .A(_05068_),
    .B(_05070_),
    .Y(_05071_)
  );
  NAND _13356_ (
    .A(_05058_),
    .B(_05071_),
    .Y(_00076_)
  );
  NAND _13357_ (
    .A(\memory[18][5] ),
    .B(_05361_),
    .Y(_05072_)
  );
  OR _13358_ (
    .A(\memory[18][5] ),
    .B(_01501_),
    .Y(_05073_)
  );
  OR _13359_ (
    .A(\data_i[29] ),
    .B(_01502_),
    .Y(_05074_)
  );
  NAND _13360_ (
    .A(_05073_),
    .B(_05074_),
    .Y(_05075_)
  );
  NAND _13361_ (
    .A(_01568_),
    .B(_05075_),
    .Y(_05076_)
  );
  OR _13362_ (
    .A(\data_i[21] ),
    .B(_01568_),
    .Y(_05077_)
  );
  AND _13363_ (
    .A(_05076_),
    .B(_05077_),
    .Y(_05078_)
  );
  NAND _13364_ (
    .A(\data_i[13] ),
    .B(_01479_),
    .Y(_05079_)
  );
  AND _13365_ (
    .A(_01583_),
    .B(_05079_),
    .Y(_05080_)
  );
  NAND _13366_ (
    .A(_01480_),
    .B(_05078_),
    .Y(_05081_)
  );
  NAND _13367_ (
    .A(_05080_),
    .B(_05081_),
    .Y(_05082_)
  );
  OR _13368_ (
    .A(\data_i[5] ),
    .B(_01583_),
    .Y(_05083_)
  );
  AND _13369_ (
    .A(MemWrite_i),
    .B(_05083_),
    .Y(_05084_)
  );
  NAND _13370_ (
    .A(_05082_),
    .B(_05084_),
    .Y(_05085_)
  );
  NAND _13371_ (
    .A(_05072_),
    .B(_05085_),
    .Y(_00077_)
  );
  OR _13372_ (
    .A(\memory[18][6] ),
    .B(MemWrite_i),
    .Y(_05086_)
  );
  NAND _13373_ (
    .A(\data_i[30] ),
    .B(_01501_),
    .Y(_05087_)
  );
  NAND _13374_ (
    .A(\memory[18][6] ),
    .B(_01502_),
    .Y(_05088_)
  );
  NAND _13375_ (
    .A(_05087_),
    .B(_05088_),
    .Y(_05089_)
  );
  NAND _13376_ (
    .A(_01568_),
    .B(_05089_),
    .Y(_05090_)
  );
  NAND _13377_ (
    .A(\data_i[22] ),
    .B(_01567_),
    .Y(_05091_)
  );
  AND _13378_ (
    .A(_01480_),
    .B(_05091_),
    .Y(_05092_)
  );
  NAND _13379_ (
    .A(_05090_),
    .B(_05092_),
    .Y(_05093_)
  );
  OR _13380_ (
    .A(\data_i[14] ),
    .B(_01480_),
    .Y(_05094_)
  );
  AND _13381_ (
    .A(_01583_),
    .B(_05094_),
    .Y(_05095_)
  );
  NAND _13382_ (
    .A(_05093_),
    .B(_05095_),
    .Y(_05096_)
  );
  NAND _13383_ (
    .A(\data_i[6] ),
    .B(_01582_),
    .Y(_05097_)
  );
  AND _13384_ (
    .A(MemWrite_i),
    .B(_05097_),
    .Y(_05098_)
  );
  NAND _13385_ (
    .A(_05096_),
    .B(_05098_),
    .Y(_05099_)
  );
  AND _13386_ (
    .A(_05086_),
    .B(_05099_),
    .Y(_00078_)
  );
  OR _13387_ (
    .A(\memory[18][7] ),
    .B(MemWrite_i),
    .Y(_05100_)
  );
  NAND _13388_ (
    .A(\data_i[31] ),
    .B(_01501_),
    .Y(_05101_)
  );
  NAND _13389_ (
    .A(\memory[18][7] ),
    .B(_01502_),
    .Y(_05102_)
  );
  NAND _13390_ (
    .A(_05101_),
    .B(_05102_),
    .Y(_05103_)
  );
  NAND _13391_ (
    .A(_01568_),
    .B(_05103_),
    .Y(_05104_)
  );
  NAND _13392_ (
    .A(\data_i[23] ),
    .B(_01567_),
    .Y(_05105_)
  );
  AND _13393_ (
    .A(_01480_),
    .B(_05105_),
    .Y(_05106_)
  );
  NAND _13394_ (
    .A(_05104_),
    .B(_05106_),
    .Y(_05107_)
  );
  OR _13395_ (
    .A(\data_i[15] ),
    .B(_01480_),
    .Y(_05108_)
  );
  AND _13396_ (
    .A(_01583_),
    .B(_05108_),
    .Y(_05109_)
  );
  NAND _13397_ (
    .A(_05107_),
    .B(_05109_),
    .Y(_05110_)
  );
  NAND _13398_ (
    .A(\data_i[7] ),
    .B(_01582_),
    .Y(_05111_)
  );
  AND _13399_ (
    .A(MemWrite_i),
    .B(_05111_),
    .Y(_05112_)
  );
  NAND _13400_ (
    .A(_05110_),
    .B(_05112_),
    .Y(_05113_)
  );
  AND _13401_ (
    .A(_05100_),
    .B(_05113_),
    .Y(_00079_)
  );
  NAND _13402_ (
    .A(\memory[17][0] ),
    .B(_05361_),
    .Y(_05114_)
  );
  OR _13403_ (
    .A(\memory[17][0] ),
    .B(_01543_),
    .Y(_05115_)
  );
  OR _13404_ (
    .A(\data_i[24] ),
    .B(_01544_),
    .Y(_05116_)
  );
  NAND _13405_ (
    .A(_05115_),
    .B(_05116_),
    .Y(_05117_)
  );
  NAND _13406_ (
    .A(_01502_),
    .B(_05117_),
    .Y(_05118_)
  );
  OR _13407_ (
    .A(\data_i[16] ),
    .B(_01502_),
    .Y(_05119_)
  );
  AND _13408_ (
    .A(_05118_),
    .B(_05119_),
    .Y(_05120_)
  );
  NAND _13409_ (
    .A(\data_i[8] ),
    .B(_01567_),
    .Y(_05121_)
  );
  AND _13410_ (
    .A(_01480_),
    .B(_05121_),
    .Y(_05122_)
  );
  NAND _13411_ (
    .A(_01568_),
    .B(_05120_),
    .Y(_05123_)
  );
  NAND _13412_ (
    .A(_05122_),
    .B(_05123_),
    .Y(_05124_)
  );
  OR _13413_ (
    .A(\data_i[0] ),
    .B(_01480_),
    .Y(_05125_)
  );
  AND _13414_ (
    .A(MemWrite_i),
    .B(_05125_),
    .Y(_05126_)
  );
  NAND _13415_ (
    .A(_05124_),
    .B(_05126_),
    .Y(_05127_)
  );
  NAND _13416_ (
    .A(_05114_),
    .B(_05127_),
    .Y(_00064_)
  );
  NAND _13417_ (
    .A(\memory[17][1] ),
    .B(_05361_),
    .Y(_05128_)
  );
  OR _13418_ (
    .A(\memory[17][1] ),
    .B(_01543_),
    .Y(_05129_)
  );
  OR _13419_ (
    .A(\data_i[25] ),
    .B(_01544_),
    .Y(_05130_)
  );
  NAND _13420_ (
    .A(_05129_),
    .B(_05130_),
    .Y(_05131_)
  );
  NAND _13421_ (
    .A(_01502_),
    .B(_05131_),
    .Y(_05132_)
  );
  OR _13422_ (
    .A(\data_i[17] ),
    .B(_01502_),
    .Y(_05133_)
  );
  AND _13423_ (
    .A(_05132_),
    .B(_05133_),
    .Y(_05134_)
  );
  NAND _13424_ (
    .A(\data_i[9] ),
    .B(_01567_),
    .Y(_05135_)
  );
  AND _13425_ (
    .A(_01480_),
    .B(_05135_),
    .Y(_05136_)
  );
  NAND _13426_ (
    .A(_01568_),
    .B(_05134_),
    .Y(_05137_)
  );
  NAND _13427_ (
    .A(_05136_),
    .B(_05137_),
    .Y(_05138_)
  );
  OR _13428_ (
    .A(\data_i[1] ),
    .B(_01480_),
    .Y(_05139_)
  );
  AND _13429_ (
    .A(MemWrite_i),
    .B(_05139_),
    .Y(_05140_)
  );
  NAND _13430_ (
    .A(_05138_),
    .B(_05140_),
    .Y(_05141_)
  );
  NAND _13431_ (
    .A(_05128_),
    .B(_05141_),
    .Y(_00065_)
  );
  NAND _13432_ (
    .A(\memory[17][2] ),
    .B(_05361_),
    .Y(_05142_)
  );
  OR _13433_ (
    .A(\memory[17][2] ),
    .B(_01543_),
    .Y(_05143_)
  );
  OR _13434_ (
    .A(\data_i[26] ),
    .B(_01544_),
    .Y(_05144_)
  );
  NAND _13435_ (
    .A(_05143_),
    .B(_05144_),
    .Y(_05145_)
  );
  NAND _13436_ (
    .A(_01502_),
    .B(_05145_),
    .Y(_05146_)
  );
  OR _13437_ (
    .A(\data_i[18] ),
    .B(_01502_),
    .Y(_05147_)
  );
  AND _13438_ (
    .A(_05146_),
    .B(_05147_),
    .Y(_05148_)
  );
  NAND _13439_ (
    .A(\data_i[10] ),
    .B(_01567_),
    .Y(_05149_)
  );
  AND _13440_ (
    .A(_01480_),
    .B(_05149_),
    .Y(_05150_)
  );
  NAND _13441_ (
    .A(_01568_),
    .B(_05148_),
    .Y(_05151_)
  );
  NAND _13442_ (
    .A(_05150_),
    .B(_05151_),
    .Y(_05152_)
  );
  OR _13443_ (
    .A(\data_i[2] ),
    .B(_01480_),
    .Y(_05153_)
  );
  AND _13444_ (
    .A(MemWrite_i),
    .B(_05153_),
    .Y(_05154_)
  );
  NAND _13445_ (
    .A(_05152_),
    .B(_05154_),
    .Y(_05155_)
  );
  NAND _13446_ (
    .A(_05142_),
    .B(_05155_),
    .Y(_00066_)
  );
  NAND _13447_ (
    .A(\memory[17][3] ),
    .B(_05361_),
    .Y(_05156_)
  );
  OR _13448_ (
    .A(\memory[17][3] ),
    .B(_01543_),
    .Y(_05157_)
  );
  OR _13449_ (
    .A(\data_i[27] ),
    .B(_01544_),
    .Y(_05158_)
  );
  NAND _13450_ (
    .A(_05157_),
    .B(_05158_),
    .Y(_05159_)
  );
  NAND _13451_ (
    .A(_01502_),
    .B(_05159_),
    .Y(_05160_)
  );
  OR _13452_ (
    .A(\data_i[19] ),
    .B(_01502_),
    .Y(_05161_)
  );
  AND _13453_ (
    .A(_05160_),
    .B(_05161_),
    .Y(_05162_)
  );
  NAND _13454_ (
    .A(\data_i[11] ),
    .B(_01567_),
    .Y(_05163_)
  );
  AND _13455_ (
    .A(_01480_),
    .B(_05163_),
    .Y(_05164_)
  );
  NAND _13456_ (
    .A(_01568_),
    .B(_05162_),
    .Y(_05165_)
  );
  NAND _13457_ (
    .A(_05164_),
    .B(_05165_),
    .Y(_05166_)
  );
  OR _13458_ (
    .A(\data_i[3] ),
    .B(_01480_),
    .Y(_05167_)
  );
  AND _13459_ (
    .A(MemWrite_i),
    .B(_05167_),
    .Y(_05168_)
  );
  NAND _13460_ (
    .A(_05166_),
    .B(_05168_),
    .Y(_05169_)
  );
  NAND _13461_ (
    .A(_05156_),
    .B(_05169_),
    .Y(_00067_)
  );
  NAND _13462_ (
    .A(\memory[17][4] ),
    .B(_05361_),
    .Y(_05170_)
  );
  OR _13463_ (
    .A(\memory[17][4] ),
    .B(_01543_),
    .Y(_05171_)
  );
  OR _13464_ (
    .A(\data_i[28] ),
    .B(_01544_),
    .Y(_05172_)
  );
  NAND _13465_ (
    .A(_05171_),
    .B(_05172_),
    .Y(_05173_)
  );
  NAND _13466_ (
    .A(_01502_),
    .B(_05173_),
    .Y(_05174_)
  );
  OR _13467_ (
    .A(\data_i[20] ),
    .B(_01502_),
    .Y(_05175_)
  );
  AND _13468_ (
    .A(_05174_),
    .B(_05175_),
    .Y(_05176_)
  );
  NAND _13469_ (
    .A(\data_i[12] ),
    .B(_01567_),
    .Y(_05177_)
  );
  AND _13470_ (
    .A(_01480_),
    .B(_05177_),
    .Y(_05178_)
  );
  NAND _13471_ (
    .A(_01568_),
    .B(_05176_),
    .Y(_05179_)
  );
  NAND _13472_ (
    .A(_05178_),
    .B(_05179_),
    .Y(_05180_)
  );
  OR _13473_ (
    .A(\data_i[4] ),
    .B(_01480_),
    .Y(_05181_)
  );
  AND _13474_ (
    .A(MemWrite_i),
    .B(_05181_),
    .Y(_05182_)
  );
  NAND _13475_ (
    .A(_05180_),
    .B(_05182_),
    .Y(_05183_)
  );
  NAND _13476_ (
    .A(_05170_),
    .B(_05183_),
    .Y(_00068_)
  );
  NAND _13477_ (
    .A(\memory[17][5] ),
    .B(_05361_),
    .Y(_05184_)
  );
  OR _13478_ (
    .A(\memory[17][5] ),
    .B(_01543_),
    .Y(_05185_)
  );
  OR _13479_ (
    .A(\data_i[29] ),
    .B(_01544_),
    .Y(_05186_)
  );
  NAND _13480_ (
    .A(_05185_),
    .B(_05186_),
    .Y(_05187_)
  );
  NAND _13481_ (
    .A(_01502_),
    .B(_05187_),
    .Y(_05188_)
  );
  OR _13482_ (
    .A(\data_i[21] ),
    .B(_01502_),
    .Y(_05189_)
  );
  AND _13483_ (
    .A(_05188_),
    .B(_05189_),
    .Y(_05190_)
  );
  NAND _13484_ (
    .A(\data_i[13] ),
    .B(_01567_),
    .Y(_05191_)
  );
  AND _13485_ (
    .A(_01480_),
    .B(_05191_),
    .Y(_05192_)
  );
  NAND _13486_ (
    .A(_01568_),
    .B(_05190_),
    .Y(_05193_)
  );
  NAND _13487_ (
    .A(_05192_),
    .B(_05193_),
    .Y(_05194_)
  );
  OR _13488_ (
    .A(\data_i[5] ),
    .B(_01480_),
    .Y(_05195_)
  );
  AND _13489_ (
    .A(MemWrite_i),
    .B(_05195_),
    .Y(_05196_)
  );
  NAND _13490_ (
    .A(_05194_),
    .B(_05196_),
    .Y(_05197_)
  );
  NAND _13491_ (
    .A(_05184_),
    .B(_05197_),
    .Y(_00069_)
  );
  NAND _13492_ (
    .A(\memory[17][6] ),
    .B(_05361_),
    .Y(_05198_)
  );
  OR _13493_ (
    .A(\memory[17][6] ),
    .B(_01543_),
    .Y(_05199_)
  );
  OR _13494_ (
    .A(\data_i[30] ),
    .B(_01544_),
    .Y(_05200_)
  );
  NAND _13495_ (
    .A(_05199_),
    .B(_05200_),
    .Y(_05201_)
  );
  NAND _13496_ (
    .A(_01502_),
    .B(_05201_),
    .Y(_05202_)
  );
  OR _13497_ (
    .A(\data_i[22] ),
    .B(_01502_),
    .Y(_05203_)
  );
  AND _13498_ (
    .A(_05202_),
    .B(_05203_),
    .Y(_05204_)
  );
  NAND _13499_ (
    .A(\data_i[14] ),
    .B(_01567_),
    .Y(_05205_)
  );
  AND _13500_ (
    .A(_01480_),
    .B(_05205_),
    .Y(_05206_)
  );
  NAND _13501_ (
    .A(_01568_),
    .B(_05204_),
    .Y(_05207_)
  );
  NAND _13502_ (
    .A(_05206_),
    .B(_05207_),
    .Y(_05208_)
  );
  OR _13503_ (
    .A(\data_i[6] ),
    .B(_01480_),
    .Y(_05209_)
  );
  AND _13504_ (
    .A(MemWrite_i),
    .B(_05209_),
    .Y(_05210_)
  );
  NAND _13505_ (
    .A(_05208_),
    .B(_05210_),
    .Y(_05211_)
  );
  NAND _13506_ (
    .A(_05198_),
    .B(_05211_),
    .Y(_00070_)
  );
  NAND _13507_ (
    .A(\memory[17][7] ),
    .B(_05361_),
    .Y(_05212_)
  );
  OR _13508_ (
    .A(\memory[17][7] ),
    .B(_01543_),
    .Y(_05213_)
  );
  OR _13509_ (
    .A(\data_i[31] ),
    .B(_01544_),
    .Y(_05214_)
  );
  NAND _13510_ (
    .A(_05213_),
    .B(_05214_),
    .Y(_05215_)
  );
  NAND _13511_ (
    .A(_01502_),
    .B(_05215_),
    .Y(_05216_)
  );
  OR _13512_ (
    .A(\data_i[23] ),
    .B(_01502_),
    .Y(_05217_)
  );
  AND _13513_ (
    .A(_05216_),
    .B(_05217_),
    .Y(_05218_)
  );
  NAND _13514_ (
    .A(\data_i[15] ),
    .B(_01567_),
    .Y(_05219_)
  );
  AND _13515_ (
    .A(_01480_),
    .B(_05219_),
    .Y(_05220_)
  );
  NAND _13516_ (
    .A(_01568_),
    .B(_05218_),
    .Y(_05221_)
  );
  NAND _13517_ (
    .A(_05220_),
    .B(_05221_),
    .Y(_05222_)
  );
  OR _13518_ (
    .A(\data_i[7] ),
    .B(_01480_),
    .Y(_05223_)
  );
  AND _13519_ (
    .A(MemWrite_i),
    .B(_05223_),
    .Y(_05224_)
  );
  NAND _13520_ (
    .A(_05222_),
    .B(_05224_),
    .Y(_05225_)
  );
  NAND _13521_ (
    .A(_05212_),
    .B(_05225_),
    .Y(_00071_)
  );
  NAND _13522_ (
    .A(\memory[16][0] ),
    .B(_05361_),
    .Y(_05226_)
  );
  OR _13523_ (
    .A(\memory[16][0] ),
    .B(_01520_),
    .Y(_05227_)
  );
  OR _13524_ (
    .A(\data_i[24] ),
    .B(_01521_),
    .Y(_05228_)
  );
  NAND _13525_ (
    .A(_05227_),
    .B(_05228_),
    .Y(_05229_)
  );
  NAND _13526_ (
    .A(_01544_),
    .B(_05229_),
    .Y(_05230_)
  );
  OR _13527_ (
    .A(\data_i[16] ),
    .B(_01544_),
    .Y(_05231_)
  );
  AND _13528_ (
    .A(_05230_),
    .B(_05231_),
    .Y(_05232_)
  );
  NAND _13529_ (
    .A(\data_i[8] ),
    .B(_01501_),
    .Y(_05233_)
  );
  AND _13530_ (
    .A(_01568_),
    .B(_05233_),
    .Y(_05234_)
  );
  NAND _13531_ (
    .A(_01502_),
    .B(_05232_),
    .Y(_05235_)
  );
  NAND _13532_ (
    .A(_05234_),
    .B(_05235_),
    .Y(_05236_)
  );
  OR _13533_ (
    .A(\data_i[0] ),
    .B(_01568_),
    .Y(_05237_)
  );
  AND _13534_ (
    .A(MemWrite_i),
    .B(_05237_),
    .Y(_05238_)
  );
  NAND _13535_ (
    .A(_05236_),
    .B(_05238_),
    .Y(_05239_)
  );
  NAND _13536_ (
    .A(_05226_),
    .B(_05239_),
    .Y(_00056_)
  );
  NAND _13537_ (
    .A(\memory[16][1] ),
    .B(_05361_),
    .Y(_05240_)
  );
  OR _13538_ (
    .A(\memory[16][1] ),
    .B(_01520_),
    .Y(_05241_)
  );
  OR _13539_ (
    .A(\data_i[25] ),
    .B(_01521_),
    .Y(_05242_)
  );
  NAND _13540_ (
    .A(_05241_),
    .B(_05242_),
    .Y(_05243_)
  );
  NAND _13541_ (
    .A(_01544_),
    .B(_05243_),
    .Y(_05244_)
  );
  OR _13542_ (
    .A(\data_i[17] ),
    .B(_01544_),
    .Y(_05245_)
  );
  AND _13543_ (
    .A(_05244_),
    .B(_05245_),
    .Y(_05246_)
  );
  NAND _13544_ (
    .A(\data_i[9] ),
    .B(_01501_),
    .Y(_05247_)
  );
  AND _13545_ (
    .A(_01568_),
    .B(_05247_),
    .Y(_05248_)
  );
  NAND _13546_ (
    .A(_01502_),
    .B(_05246_),
    .Y(_05249_)
  );
  NAND _13547_ (
    .A(_05248_),
    .B(_05249_),
    .Y(_05250_)
  );
  OR _13548_ (
    .A(\data_i[1] ),
    .B(_01568_),
    .Y(_05251_)
  );
  AND _13549_ (
    .A(MemWrite_i),
    .B(_05251_),
    .Y(_05252_)
  );
  NAND _13550_ (
    .A(_05250_),
    .B(_05252_),
    .Y(_05253_)
  );
  NAND _13551_ (
    .A(_05240_),
    .B(_05253_),
    .Y(_00057_)
  );
  NAND _13552_ (
    .A(\memory[16][2] ),
    .B(_05361_),
    .Y(_05254_)
  );
  OR _13553_ (
    .A(\memory[16][2] ),
    .B(_01520_),
    .Y(_05255_)
  );
  OR _13554_ (
    .A(\data_i[26] ),
    .B(_01521_),
    .Y(_05256_)
  );
  NAND _13555_ (
    .A(_05255_),
    .B(_05256_),
    .Y(_05257_)
  );
  NAND _13556_ (
    .A(_01544_),
    .B(_05257_),
    .Y(_05258_)
  );
  OR _13557_ (
    .A(\data_i[18] ),
    .B(_01544_),
    .Y(_05259_)
  );
  AND _13558_ (
    .A(_05258_),
    .B(_05259_),
    .Y(_05260_)
  );
  NAND _13559_ (
    .A(\data_i[10] ),
    .B(_01501_),
    .Y(_05261_)
  );
  AND _13560_ (
    .A(_01568_),
    .B(_05261_),
    .Y(_05262_)
  );
  NAND _13561_ (
    .A(_01502_),
    .B(_05260_),
    .Y(_05263_)
  );
  NAND _13562_ (
    .A(_05262_),
    .B(_05263_),
    .Y(_05264_)
  );
  OR _13563_ (
    .A(\data_i[2] ),
    .B(_01568_),
    .Y(_05265_)
  );
  AND _13564_ (
    .A(MemWrite_i),
    .B(_05265_),
    .Y(_05266_)
  );
  NAND _13565_ (
    .A(_05264_),
    .B(_05266_),
    .Y(_05267_)
  );
  NAND _13566_ (
    .A(_05254_),
    .B(_05267_),
    .Y(_00058_)
  );
  NAND _13567_ (
    .A(\memory[16][3] ),
    .B(_05361_),
    .Y(_05268_)
  );
  OR _13568_ (
    .A(\memory[16][3] ),
    .B(_01520_),
    .Y(_05269_)
  );
  OR _13569_ (
    .A(\data_i[27] ),
    .B(_01521_),
    .Y(_05270_)
  );
  NAND _13570_ (
    .A(_05269_),
    .B(_05270_),
    .Y(_05271_)
  );
  NAND _13571_ (
    .A(_01544_),
    .B(_05271_),
    .Y(_05272_)
  );
  OR _13572_ (
    .A(\data_i[19] ),
    .B(_01544_),
    .Y(_05273_)
  );
  AND _13573_ (
    .A(_05272_),
    .B(_05273_),
    .Y(_05274_)
  );
  NAND _13574_ (
    .A(\data_i[11] ),
    .B(_01501_),
    .Y(_05275_)
  );
  AND _13575_ (
    .A(_01568_),
    .B(_05275_),
    .Y(_05276_)
  );
  NAND _13576_ (
    .A(_01502_),
    .B(_05274_),
    .Y(_05277_)
  );
  NAND _13577_ (
    .A(_05276_),
    .B(_05277_),
    .Y(_05278_)
  );
  OR _13578_ (
    .A(\data_i[3] ),
    .B(_01568_),
    .Y(_05279_)
  );
  AND _13579_ (
    .A(MemWrite_i),
    .B(_05279_),
    .Y(_05280_)
  );
  NAND _13580_ (
    .A(_05278_),
    .B(_05280_),
    .Y(_05281_)
  );
  NAND _13581_ (
    .A(_05268_),
    .B(_05281_),
    .Y(_00059_)
  );
  NAND _13582_ (
    .A(\memory[16][4] ),
    .B(_05361_),
    .Y(_05282_)
  );
  OR _13583_ (
    .A(\memory[16][4] ),
    .B(_01520_),
    .Y(_05283_)
  );
  OR _13584_ (
    .A(\data_i[28] ),
    .B(_01521_),
    .Y(_05284_)
  );
  NAND _13585_ (
    .A(_05283_),
    .B(_05284_),
    .Y(_05285_)
  );
  NAND _13586_ (
    .A(_01544_),
    .B(_05285_),
    .Y(_05286_)
  );
  OR _13587_ (
    .A(\data_i[20] ),
    .B(_01544_),
    .Y(_05287_)
  );
  AND _13588_ (
    .A(_05286_),
    .B(_05287_),
    .Y(_05288_)
  );
  NAND _13589_ (
    .A(\data_i[12] ),
    .B(_01501_),
    .Y(_05289_)
  );
  AND _13590_ (
    .A(_01568_),
    .B(_05289_),
    .Y(_05290_)
  );
  NAND _13591_ (
    .A(_01502_),
    .B(_05288_),
    .Y(_05291_)
  );
  NAND _13592_ (
    .A(_05290_),
    .B(_05291_),
    .Y(_05292_)
  );
  OR _13593_ (
    .A(\data_i[4] ),
    .B(_01568_),
    .Y(_05293_)
  );
  AND _13594_ (
    .A(MemWrite_i),
    .B(_05293_),
    .Y(_05294_)
  );
  NAND _13595_ (
    .A(_05292_),
    .B(_05294_),
    .Y(_05295_)
  );
  NAND _13596_ (
    .A(_05282_),
    .B(_05295_),
    .Y(_00060_)
  );
  NAND _13597_ (
    .A(\memory[16][5] ),
    .B(_05361_),
    .Y(_05296_)
  );
  OR _13598_ (
    .A(\memory[16][5] ),
    .B(_01520_),
    .Y(_05297_)
  );
  OR _13599_ (
    .A(\data_i[29] ),
    .B(_01521_),
    .Y(_05298_)
  );
  NAND _13600_ (
    .A(_05297_),
    .B(_05298_),
    .Y(_05300_)
  );
  NAND _13601_ (
    .A(_01544_),
    .B(_05300_),
    .Y(_05301_)
  );
  OR _13602_ (
    .A(\data_i[21] ),
    .B(_01544_),
    .Y(_05302_)
  );
  AND _13603_ (
    .A(_05301_),
    .B(_05302_),
    .Y(_05303_)
  );
  NAND _13604_ (
    .A(\data_i[13] ),
    .B(_01501_),
    .Y(_05304_)
  );
  AND _13605_ (
    .A(_01568_),
    .B(_05304_),
    .Y(_05305_)
  );
  NAND _13606_ (
    .A(_01502_),
    .B(_05303_),
    .Y(_05306_)
  );
  NAND _13607_ (
    .A(_05305_),
    .B(_05306_),
    .Y(_05307_)
  );
  OR _13608_ (
    .A(\data_i[5] ),
    .B(_01568_),
    .Y(_05308_)
  );
  AND _13609_ (
    .A(MemWrite_i),
    .B(_05308_),
    .Y(_05309_)
  );
  NAND _13610_ (
    .A(_05307_),
    .B(_05309_),
    .Y(_05311_)
  );
  NAND _13611_ (
    .A(_05296_),
    .B(_05311_),
    .Y(_00061_)
  );
  NAND _13612_ (
    .A(\memory[16][6] ),
    .B(_05361_),
    .Y(_05312_)
  );
  OR _13613_ (
    .A(\memory[16][6] ),
    .B(_01520_),
    .Y(_05313_)
  );
  OR _13614_ (
    .A(\data_i[30] ),
    .B(_01521_),
    .Y(_05314_)
  );
  NAND _13615_ (
    .A(_05313_),
    .B(_05314_),
    .Y(_05315_)
  );
  NAND _13616_ (
    .A(_01544_),
    .B(_05315_),
    .Y(_05316_)
  );
  OR _13617_ (
    .A(\data_i[22] ),
    .B(_01544_),
    .Y(_05317_)
  );
  AND _13618_ (
    .A(_05316_),
    .B(_05317_),
    .Y(_05318_)
  );
  NAND _13619_ (
    .A(\data_i[14] ),
    .B(_01501_),
    .Y(_05319_)
  );
  AND _13620_ (
    .A(_01568_),
    .B(_05319_),
    .Y(_05321_)
  );
  NAND _13621_ (
    .A(_01502_),
    .B(_05318_),
    .Y(_05322_)
  );
  NAND _13622_ (
    .A(_05321_),
    .B(_05322_),
    .Y(_05323_)
  );
  OR _13623_ (
    .A(\data_i[6] ),
    .B(_01568_),
    .Y(_05324_)
  );
  AND _13624_ (
    .A(MemWrite_i),
    .B(_05324_),
    .Y(_05325_)
  );
  NAND _13625_ (
    .A(_05323_),
    .B(_05325_),
    .Y(_05326_)
  );
  NAND _13626_ (
    .A(_05312_),
    .B(_05326_),
    .Y(_00062_)
  );
  NAND _13627_ (
    .A(\memory[16][7] ),
    .B(_05361_),
    .Y(_05327_)
  );
  OR _13628_ (
    .A(\memory[16][7] ),
    .B(_01520_),
    .Y(_05328_)
  );
  OR _13629_ (
    .A(\data_i[31] ),
    .B(_01521_),
    .Y(_05329_)
  );
  NAND _13630_ (
    .A(_05328_),
    .B(_05329_),
    .Y(_05331_)
  );
  NAND _13631_ (
    .A(_01544_),
    .B(_05331_),
    .Y(_05332_)
  );
  OR _13632_ (
    .A(\data_i[23] ),
    .B(_01544_),
    .Y(_05333_)
  );
  AND _13633_ (
    .A(_05332_),
    .B(_05333_),
    .Y(_05334_)
  );
  NAND _13634_ (
    .A(\data_i[15] ),
    .B(_01501_),
    .Y(_05335_)
  );
  AND _13635_ (
    .A(_01568_),
    .B(_05335_),
    .Y(_05336_)
  );
  NAND _13636_ (
    .A(_01502_),
    .B(_05334_),
    .Y(_05337_)
  );
  NAND _13637_ (
    .A(_05336_),
    .B(_05337_),
    .Y(_05338_)
  );
  OR _13638_ (
    .A(\data_i[7] ),
    .B(_01568_),
    .Y(_05339_)
  );
  AND _13639_ (
    .A(MemWrite_i),
    .B(_05339_),
    .Y(_05340_)
  );
  NAND _13640_ (
    .A(_05338_),
    .B(_05340_),
    .Y(_05342_)
  );
  NAND _13641_ (
    .A(_05327_),
    .B(_05342_),
    .Y(_00063_)
  );
  NAND _13642_ (
    .A(\memory[15][0] ),
    .B(_05361_),
    .Y(_05343_)
  );
  OR _13643_ (
    .A(\memory[15][0] ),
    .B(_01458_),
    .Y(_05344_)
  );
  OR _13644_ (
    .A(\data_i[24] ),
    .B(_01459_),
    .Y(_05345_)
  );
  NAND _13645_ (
    .A(_05344_),
    .B(_05345_),
    .Y(_05346_)
  );
  NAND _13646_ (
    .A(_01521_),
    .B(_05346_),
    .Y(_05347_)
  );
  OR _13647_ (
    .A(\data_i[16] ),
    .B(_01521_),
    .Y(_05348_)
  );
  AND _13648_ (
    .A(_05347_),
    .B(_05348_),
    .Y(_05349_)
  );
  NAND _13649_ (
    .A(\data_i[8] ),
    .B(_01543_),
    .Y(_05350_)
  );
  AND _13650_ (
    .A(_01502_),
    .B(_05350_),
    .Y(_05352_)
  );
  NAND _13651_ (
    .A(_01544_),
    .B(_05349_),
    .Y(_05353_)
  );
  NAND _13652_ (
    .A(_05352_),
    .B(_05353_),
    .Y(_05354_)
  );
  OR _13653_ (
    .A(\data_i[0] ),
    .B(_01502_),
    .Y(_05355_)
  );
  AND _13654_ (
    .A(MemWrite_i),
    .B(_05355_),
    .Y(_05356_)
  );
  NAND _13655_ (
    .A(_05354_),
    .B(_05356_),
    .Y(_05357_)
  );
  NAND _13656_ (
    .A(_05343_),
    .B(_05357_),
    .Y(_00048_)
  );
  NAND _13657_ (
    .A(\memory[15][1] ),
    .B(_05361_),
    .Y(_05358_)
  );
  OR _13658_ (
    .A(\memory[15][1] ),
    .B(_01458_),
    .Y(_05359_)
  );
  OR _13659_ (
    .A(\data_i[25] ),
    .B(_01459_),
    .Y(_05360_)
  );
  NAND _13660_ (
    .A(_05359_),
    .B(_05360_),
    .Y(_05362_)
  );
  NAND _13661_ (
    .A(_01521_),
    .B(_05362_),
    .Y(_05363_)
  );
  OR _13662_ (
    .A(\data_i[17] ),
    .B(_01521_),
    .Y(_05364_)
  );
  AND _13663_ (
    .A(_05363_),
    .B(_05364_),
    .Y(_05365_)
  );
  NAND _13664_ (
    .A(\data_i[9] ),
    .B(_01543_),
    .Y(_05366_)
  );
  AND _13665_ (
    .A(_01502_),
    .B(_05366_),
    .Y(_05367_)
  );
  NAND _13666_ (
    .A(_01544_),
    .B(_05365_),
    .Y(_05368_)
  );
  NAND _13667_ (
    .A(_05367_),
    .B(_05368_),
    .Y(_05369_)
  );
  OR _13668_ (
    .A(\data_i[1] ),
    .B(_01502_),
    .Y(_05370_)
  );
  AND _13669_ (
    .A(MemWrite_i),
    .B(_05370_),
    .Y(_05371_)
  );
  NAND _13670_ (
    .A(_05369_),
    .B(_05371_),
    .Y(_05373_)
  );
  NAND _13671_ (
    .A(_05358_),
    .B(_05373_),
    .Y(_00049_)
  );
  NAND _13672_ (
    .A(\memory[15][2] ),
    .B(_05361_),
    .Y(_05374_)
  );
  OR _13673_ (
    .A(\memory[15][2] ),
    .B(_01458_),
    .Y(_05375_)
  );
  OR _13674_ (
    .A(\data_i[26] ),
    .B(_01459_),
    .Y(_05376_)
  );
  NAND _13675_ (
    .A(_05375_),
    .B(_05376_),
    .Y(_05377_)
  );
  NAND _13676_ (
    .A(_01521_),
    .B(_05377_),
    .Y(_05378_)
  );
  OR _13677_ (
    .A(\data_i[18] ),
    .B(_01521_),
    .Y(_05379_)
  );
  AND _13678_ (
    .A(_05378_),
    .B(_05379_),
    .Y(_05380_)
  );
  NAND _13679_ (
    .A(\data_i[10] ),
    .B(_01543_),
    .Y(_05381_)
  );
  AND _13680_ (
    .A(_01502_),
    .B(_05381_),
    .Y(_05383_)
  );
  NAND _13681_ (
    .A(_01544_),
    .B(_05380_),
    .Y(_05384_)
  );
  NAND _13682_ (
    .A(_05383_),
    .B(_05384_),
    .Y(_05385_)
  );
  OR _13683_ (
    .A(\data_i[2] ),
    .B(_01502_),
    .Y(_05386_)
  );
  AND _13684_ (
    .A(MemWrite_i),
    .B(_05386_),
    .Y(_05387_)
  );
  NAND _13685_ (
    .A(_05385_),
    .B(_05387_),
    .Y(_05388_)
  );
  NAND _13686_ (
    .A(_05374_),
    .B(_05388_),
    .Y(_00050_)
  );
  NAND _13687_ (
    .A(\memory[15][3] ),
    .B(_05361_),
    .Y(_05389_)
  );
  OR _13688_ (
    .A(\memory[15][3] ),
    .B(_01458_),
    .Y(_05390_)
  );
  OR _13689_ (
    .A(\data_i[27] ),
    .B(_01459_),
    .Y(_05391_)
  );
  NAND _13690_ (
    .A(_05390_),
    .B(_05391_),
    .Y(_05393_)
  );
  NAND _13691_ (
    .A(_01521_),
    .B(_05393_),
    .Y(_05394_)
  );
  OR _13692_ (
    .A(\data_i[19] ),
    .B(_01521_),
    .Y(_05395_)
  );
  AND _13693_ (
    .A(_05394_),
    .B(_05395_),
    .Y(_05396_)
  );
  NAND _13694_ (
    .A(\data_i[11] ),
    .B(_01543_),
    .Y(_05397_)
  );
  AND _13695_ (
    .A(_01502_),
    .B(_05397_),
    .Y(_05398_)
  );
  NAND _13696_ (
    .A(_01544_),
    .B(_05396_),
    .Y(_05399_)
  );
  NAND _13697_ (
    .A(_05398_),
    .B(_05399_),
    .Y(_05400_)
  );
  OR _13698_ (
    .A(\data_i[3] ),
    .B(_01502_),
    .Y(_05401_)
  );
  AND _13699_ (
    .A(MemWrite_i),
    .B(_05401_),
    .Y(_05402_)
  );
  NAND _13700_ (
    .A(_05400_),
    .B(_05402_),
    .Y(_05404_)
  );
  NAND _13701_ (
    .A(_05389_),
    .B(_05404_),
    .Y(_00051_)
  );
  NAND _13702_ (
    .A(\memory[15][4] ),
    .B(_05361_),
    .Y(_05405_)
  );
  OR _13703_ (
    .A(\memory[15][4] ),
    .B(_01458_),
    .Y(_05406_)
  );
  OR _13704_ (
    .A(\data_i[28] ),
    .B(_01459_),
    .Y(_05407_)
  );
  NAND _13705_ (
    .A(_05406_),
    .B(_05407_),
    .Y(_05408_)
  );
  NAND _13706_ (
    .A(_01521_),
    .B(_05408_),
    .Y(_05409_)
  );
  OR _13707_ (
    .A(\data_i[20] ),
    .B(_01521_),
    .Y(_05410_)
  );
  AND _13708_ (
    .A(_05409_),
    .B(_05410_),
    .Y(_05411_)
  );
  NAND _13709_ (
    .A(\data_i[12] ),
    .B(_01543_),
    .Y(_05412_)
  );
  AND _13710_ (
    .A(_01502_),
    .B(_05412_),
    .Y(_05414_)
  );
  NAND _13711_ (
    .A(_01544_),
    .B(_05411_),
    .Y(_05415_)
  );
  NAND _13712_ (
    .A(_05414_),
    .B(_05415_),
    .Y(_05416_)
  );
  OR _13713_ (
    .A(\data_i[4] ),
    .B(_01502_),
    .Y(_05417_)
  );
  AND _13714_ (
    .A(MemWrite_i),
    .B(_05417_),
    .Y(_05418_)
  );
  NAND _13715_ (
    .A(_05416_),
    .B(_05418_),
    .Y(_05419_)
  );
  NAND _13716_ (
    .A(_05405_),
    .B(_05419_),
    .Y(_00052_)
  );
  NAND _13717_ (
    .A(\memory[15][5] ),
    .B(_05361_),
    .Y(_05420_)
  );
  OR _13718_ (
    .A(\memory[15][5] ),
    .B(_01458_),
    .Y(_05421_)
  );
  OR _13719_ (
    .A(\data_i[29] ),
    .B(_01459_),
    .Y(_05422_)
  );
  NAND _13720_ (
    .A(_05421_),
    .B(_05422_),
    .Y(_05424_)
  );
  NAND _13721_ (
    .A(_01521_),
    .B(_05424_),
    .Y(_05425_)
  );
  OR _13722_ (
    .A(\data_i[21] ),
    .B(_01521_),
    .Y(_05426_)
  );
  AND _13723_ (
    .A(_05425_),
    .B(_05426_),
    .Y(_05427_)
  );
  NAND _13724_ (
    .A(\data_i[13] ),
    .B(_01543_),
    .Y(_05428_)
  );
  AND _13725_ (
    .A(_01502_),
    .B(_05428_),
    .Y(_05429_)
  );
  NAND _13726_ (
    .A(_01544_),
    .B(_05427_),
    .Y(_05430_)
  );
  NAND _13727_ (
    .A(_05429_),
    .B(_05430_),
    .Y(_05431_)
  );
  OR _13728_ (
    .A(\data_i[5] ),
    .B(_01502_),
    .Y(_05432_)
  );
  AND _13729_ (
    .A(MemWrite_i),
    .B(_05432_),
    .Y(_05433_)
  );
  NAND _13730_ (
    .A(_05431_),
    .B(_05433_),
    .Y(_05435_)
  );
  NAND _13731_ (
    .A(_05420_),
    .B(_05435_),
    .Y(_00053_)
  );
  NAND _13732_ (
    .A(\memory[15][6] ),
    .B(_05361_),
    .Y(_05436_)
  );
  OR _13733_ (
    .A(\memory[15][6] ),
    .B(_01458_),
    .Y(_05437_)
  );
  OR _13734_ (
    .A(\data_i[30] ),
    .B(_01459_),
    .Y(_05438_)
  );
  NAND _13735_ (
    .A(_05437_),
    .B(_05438_),
    .Y(_05439_)
  );
  NAND _13736_ (
    .A(_01521_),
    .B(_05439_),
    .Y(_05440_)
  );
  OR _13737_ (
    .A(\data_i[22] ),
    .B(_01521_),
    .Y(_05441_)
  );
  AND _13738_ (
    .A(_05440_),
    .B(_05441_),
    .Y(_05442_)
  );
  NAND _13739_ (
    .A(\data_i[14] ),
    .B(_01543_),
    .Y(_05443_)
  );
  AND _13740_ (
    .A(_01502_),
    .B(_05443_),
    .Y(_05445_)
  );
  NAND _13741_ (
    .A(_01544_),
    .B(_05442_),
    .Y(_05446_)
  );
  NAND _13742_ (
    .A(_05445_),
    .B(_05446_),
    .Y(_05447_)
  );
  OR _13743_ (
    .A(\data_i[6] ),
    .B(_01502_),
    .Y(_05448_)
  );
  AND _13744_ (
    .A(MemWrite_i),
    .B(_05448_),
    .Y(_05449_)
  );
  NAND _13745_ (
    .A(_05447_),
    .B(_05449_),
    .Y(_05450_)
  );
  NAND _13746_ (
    .A(_05436_),
    .B(_05450_),
    .Y(_00054_)
  );
  NAND _13747_ (
    .A(\memory[15][7] ),
    .B(_05361_),
    .Y(_05451_)
  );
  OR _13748_ (
    .A(\memory[15][7] ),
    .B(_01458_),
    .Y(_05452_)
  );
  OR _13749_ (
    .A(\data_i[31] ),
    .B(_01459_),
    .Y(_05453_)
  );
  NAND _13750_ (
    .A(_05452_),
    .B(_05453_),
    .Y(_05455_)
  );
  NAND _13751_ (
    .A(_01521_),
    .B(_05455_),
    .Y(_05456_)
  );
  OR _13752_ (
    .A(\data_i[23] ),
    .B(_01521_),
    .Y(_05457_)
  );
  AND _13753_ (
    .A(_05456_),
    .B(_05457_),
    .Y(_05458_)
  );
  NAND _13754_ (
    .A(\data_i[15] ),
    .B(_01543_),
    .Y(_05459_)
  );
  AND _13755_ (
    .A(_01502_),
    .B(_05459_),
    .Y(_05460_)
  );
  NAND _13756_ (
    .A(_01544_),
    .B(_05458_),
    .Y(_05461_)
  );
  NAND _13757_ (
    .A(_05460_),
    .B(_05461_),
    .Y(_05462_)
  );
  OR _13758_ (
    .A(\data_i[7] ),
    .B(_01502_),
    .Y(_05463_)
  );
  AND _13759_ (
    .A(MemWrite_i),
    .B(_05463_),
    .Y(_05464_)
  );
  NAND _13760_ (
    .A(_05462_),
    .B(_05464_),
    .Y(_05466_)
  );
  NAND _13761_ (
    .A(_05451_),
    .B(_05466_),
    .Y(_00055_)
  );
  NAND _13762_ (
    .A(\memory[14][0] ),
    .B(_05361_),
    .Y(_05467_)
  );
  OR _13763_ (
    .A(\memory[14][0] ),
    .B(_01575_),
    .Y(_05468_)
  );
  OR _13764_ (
    .A(\data_i[24] ),
    .B(_01576_),
    .Y(_05469_)
  );
  NAND _13765_ (
    .A(_05468_),
    .B(_05469_),
    .Y(_05470_)
  );
  NAND _13766_ (
    .A(_01459_),
    .B(_05470_),
    .Y(_05471_)
  );
  OR _13767_ (
    .A(\data_i[16] ),
    .B(_01459_),
    .Y(_05472_)
  );
  AND _13768_ (
    .A(_05471_),
    .B(_05472_),
    .Y(_05473_)
  );
  NAND _13769_ (
    .A(\data_i[8] ),
    .B(_01520_),
    .Y(_05474_)
  );
  AND _13770_ (
    .A(_01544_),
    .B(_05474_),
    .Y(_05476_)
  );
  NAND _13771_ (
    .A(_01521_),
    .B(_05473_),
    .Y(_05477_)
  );
  NAND _13772_ (
    .A(_05476_),
    .B(_05477_),
    .Y(_05478_)
  );
  OR _13773_ (
    .A(\data_i[0] ),
    .B(_01544_),
    .Y(_05479_)
  );
  AND _13774_ (
    .A(MemWrite_i),
    .B(_05479_),
    .Y(_05480_)
  );
  NAND _13775_ (
    .A(_05478_),
    .B(_05480_),
    .Y(_05481_)
  );
  NAND _13776_ (
    .A(_05467_),
    .B(_05481_),
    .Y(_00040_)
  );
  NAND _13777_ (
    .A(\memory[14][1] ),
    .B(_05361_),
    .Y(_05482_)
  );
  OR _13778_ (
    .A(\memory[14][1] ),
    .B(_01575_),
    .Y(_05483_)
  );
  OR _13779_ (
    .A(\data_i[25] ),
    .B(_01576_),
    .Y(_05484_)
  );
  NAND _13780_ (
    .A(_05483_),
    .B(_05484_),
    .Y(_05486_)
  );
  NAND _13781_ (
    .A(_01459_),
    .B(_05486_),
    .Y(_05487_)
  );
  OR _13782_ (
    .A(\data_i[17] ),
    .B(_01459_),
    .Y(_05488_)
  );
  AND _13783_ (
    .A(_05487_),
    .B(_05488_),
    .Y(_05489_)
  );
  NAND _13784_ (
    .A(\data_i[9] ),
    .B(_01520_),
    .Y(_05490_)
  );
  AND _13785_ (
    .A(_01544_),
    .B(_05490_),
    .Y(_05491_)
  );
  NAND _13786_ (
    .A(_01521_),
    .B(_05489_),
    .Y(_05492_)
  );
  NAND _13787_ (
    .A(_05491_),
    .B(_05492_),
    .Y(_05493_)
  );
  OR _13788_ (
    .A(\data_i[1] ),
    .B(_01544_),
    .Y(_05494_)
  );
  AND _13789_ (
    .A(MemWrite_i),
    .B(_05494_),
    .Y(_05495_)
  );
  NAND _13790_ (
    .A(_05493_),
    .B(_05495_),
    .Y(_05497_)
  );
  NAND _13791_ (
    .A(_05482_),
    .B(_05497_),
    .Y(_00041_)
  );
  NAND _13792_ (
    .A(\memory[14][2] ),
    .B(_05361_),
    .Y(_05498_)
  );
  OR _13793_ (
    .A(\memory[14][2] ),
    .B(_01575_),
    .Y(_05499_)
  );
  OR _13794_ (
    .A(\data_i[26] ),
    .B(_01576_),
    .Y(_05500_)
  );
  NAND _13795_ (
    .A(_05499_),
    .B(_05500_),
    .Y(_05501_)
  );
  NAND _13796_ (
    .A(_01459_),
    .B(_05501_),
    .Y(_05502_)
  );
  OR _13797_ (
    .A(\data_i[18] ),
    .B(_01459_),
    .Y(_05503_)
  );
  AND _13798_ (
    .A(_05502_),
    .B(_05503_),
    .Y(_05504_)
  );
  NAND _13799_ (
    .A(\data_i[10] ),
    .B(_01520_),
    .Y(_05505_)
  );
  AND _13800_ (
    .A(_01544_),
    .B(_05505_),
    .Y(_05507_)
  );
  NAND _13801_ (
    .A(_01521_),
    .B(_05504_),
    .Y(_05508_)
  );
  NAND _13802_ (
    .A(_05507_),
    .B(_05508_),
    .Y(_05509_)
  );
  OR _13803_ (
    .A(\data_i[2] ),
    .B(_01544_),
    .Y(_05510_)
  );
  AND _13804_ (
    .A(MemWrite_i),
    .B(_05510_),
    .Y(_05511_)
  );
  NAND _13805_ (
    .A(_05509_),
    .B(_05511_),
    .Y(_05512_)
  );
  NAND _13806_ (
    .A(_05498_),
    .B(_05512_),
    .Y(_00042_)
  );
  NAND _13807_ (
    .A(\memory[14][3] ),
    .B(_05361_),
    .Y(_05513_)
  );
  OR _13808_ (
    .A(\memory[14][3] ),
    .B(_01575_),
    .Y(_05514_)
  );
  OR _13809_ (
    .A(\data_i[27] ),
    .B(_01576_),
    .Y(_05515_)
  );
  NAND _13810_ (
    .A(_05514_),
    .B(_05515_),
    .Y(_05517_)
  );
  NAND _13811_ (
    .A(_01459_),
    .B(_05517_),
    .Y(_05518_)
  );
  OR _13812_ (
    .A(\data_i[19] ),
    .B(_01459_),
    .Y(_05519_)
  );
  AND _13813_ (
    .A(_05518_),
    .B(_05519_),
    .Y(_05520_)
  );
  NAND _13814_ (
    .A(\data_i[11] ),
    .B(_01520_),
    .Y(_05521_)
  );
  AND _13815_ (
    .A(_01544_),
    .B(_05521_),
    .Y(_05522_)
  );
  NAND _13816_ (
    .A(_01521_),
    .B(_05520_),
    .Y(_05523_)
  );
  NAND _13817_ (
    .A(_05522_),
    .B(_05523_),
    .Y(_05524_)
  );
  OR _13818_ (
    .A(\data_i[3] ),
    .B(_01544_),
    .Y(_05525_)
  );
  AND _13819_ (
    .A(MemWrite_i),
    .B(_05525_),
    .Y(_05526_)
  );
  NAND _13820_ (
    .A(_05524_),
    .B(_05526_),
    .Y(_05528_)
  );
  NAND _13821_ (
    .A(_05513_),
    .B(_05528_),
    .Y(_00043_)
  );
  NAND _13822_ (
    .A(\memory[14][4] ),
    .B(_05361_),
    .Y(_05529_)
  );
  OR _13823_ (
    .A(\memory[14][4] ),
    .B(_01575_),
    .Y(_05530_)
  );
  OR _13824_ (
    .A(\data_i[28] ),
    .B(_01576_),
    .Y(_05531_)
  );
  NAND _13825_ (
    .A(_05530_),
    .B(_05531_),
    .Y(_05532_)
  );
  NAND _13826_ (
    .A(_01459_),
    .B(_05532_),
    .Y(_05533_)
  );
  OR _13827_ (
    .A(\data_i[20] ),
    .B(_01459_),
    .Y(_05534_)
  );
  AND _13828_ (
    .A(_05533_),
    .B(_05534_),
    .Y(_05535_)
  );
  NAND _13829_ (
    .A(\data_i[12] ),
    .B(_01520_),
    .Y(_05536_)
  );
  AND _13830_ (
    .A(_01544_),
    .B(_05536_),
    .Y(_05538_)
  );
  NAND _13831_ (
    .A(_01521_),
    .B(_05535_),
    .Y(_05539_)
  );
  NAND _13832_ (
    .A(_05538_),
    .B(_05539_),
    .Y(_05540_)
  );
  OR _13833_ (
    .A(\data_i[4] ),
    .B(_01544_),
    .Y(_05541_)
  );
  AND _13834_ (
    .A(MemWrite_i),
    .B(_05541_),
    .Y(_05542_)
  );
  NAND _13835_ (
    .A(_05540_),
    .B(_05542_),
    .Y(_05543_)
  );
  NAND _13836_ (
    .A(_05529_),
    .B(_05543_),
    .Y(_00044_)
  );
  NAND _13837_ (
    .A(\memory[14][5] ),
    .B(_05361_),
    .Y(_05544_)
  );
  OR _13838_ (
    .A(\memory[14][5] ),
    .B(_01575_),
    .Y(_05545_)
  );
  OR _13839_ (
    .A(\data_i[29] ),
    .B(_01576_),
    .Y(_05546_)
  );
  NAND _13840_ (
    .A(_05545_),
    .B(_05546_),
    .Y(_05548_)
  );
  NAND _13841_ (
    .A(_01459_),
    .B(_05548_),
    .Y(_05549_)
  );
  OR _13842_ (
    .A(\data_i[21] ),
    .B(_01459_),
    .Y(_05550_)
  );
  AND _13843_ (
    .A(_05549_),
    .B(_05550_),
    .Y(_05551_)
  );
  NAND _13844_ (
    .A(\data_i[13] ),
    .B(_01520_),
    .Y(_05552_)
  );
  AND _13845_ (
    .A(_01544_),
    .B(_05552_),
    .Y(_05553_)
  );
  NAND _13846_ (
    .A(_01521_),
    .B(_05551_),
    .Y(_05554_)
  );
  NAND _13847_ (
    .A(_05553_),
    .B(_05554_),
    .Y(_05555_)
  );
  OR _13848_ (
    .A(\data_i[5] ),
    .B(_01544_),
    .Y(_05556_)
  );
  AND _13849_ (
    .A(MemWrite_i),
    .B(_05556_),
    .Y(_05557_)
  );
  NAND _13850_ (
    .A(_05555_),
    .B(_05557_),
    .Y(_05559_)
  );
  NAND _13851_ (
    .A(_05544_),
    .B(_05559_),
    .Y(_00045_)
  );
  NAND _13852_ (
    .A(\memory[14][6] ),
    .B(_05361_),
    .Y(_05560_)
  );
  OR _13853_ (
    .A(\memory[14][6] ),
    .B(_01575_),
    .Y(_05561_)
  );
  OR _13854_ (
    .A(\data_i[30] ),
    .B(_01576_),
    .Y(_05562_)
  );
  NAND _13855_ (
    .A(_05561_),
    .B(_05562_),
    .Y(_05563_)
  );
  NAND _13856_ (
    .A(_01459_),
    .B(_05563_),
    .Y(_05564_)
  );
  OR _13857_ (
    .A(\data_i[22] ),
    .B(_01459_),
    .Y(_05565_)
  );
  AND _13858_ (
    .A(_05564_),
    .B(_05565_),
    .Y(_05566_)
  );
  NAND _13859_ (
    .A(\data_i[14] ),
    .B(_01520_),
    .Y(_05567_)
  );
  AND _13860_ (
    .A(_01544_),
    .B(_05567_),
    .Y(_05569_)
  );
  NAND _13861_ (
    .A(_01521_),
    .B(_05566_),
    .Y(_05570_)
  );
  NAND _13862_ (
    .A(_05569_),
    .B(_05570_),
    .Y(_05571_)
  );
  OR _13863_ (
    .A(\data_i[6] ),
    .B(_01544_),
    .Y(_05572_)
  );
  AND _13864_ (
    .A(MemWrite_i),
    .B(_05572_),
    .Y(_05573_)
  );
  NAND _13865_ (
    .A(_05571_),
    .B(_05573_),
    .Y(_05574_)
  );
  NAND _13866_ (
    .A(_05560_),
    .B(_05574_),
    .Y(_00046_)
  );
  NAND _13867_ (
    .A(\memory[14][7] ),
    .B(_05361_),
    .Y(_05575_)
  );
  OR _13868_ (
    .A(\memory[14][7] ),
    .B(_01575_),
    .Y(_05576_)
  );
  OR _13869_ (
    .A(\data_i[31] ),
    .B(_01576_),
    .Y(_05577_)
  );
  NAND _13870_ (
    .A(_05576_),
    .B(_05577_),
    .Y(_05579_)
  );
  NAND _13871_ (
    .A(_01459_),
    .B(_05579_),
    .Y(_05580_)
  );
  OR _13872_ (
    .A(\data_i[23] ),
    .B(_01459_),
    .Y(_05581_)
  );
  AND _13873_ (
    .A(_05580_),
    .B(_05581_),
    .Y(_05582_)
  );
  NAND _13874_ (
    .A(\data_i[15] ),
    .B(_01520_),
    .Y(_05583_)
  );
  AND _13875_ (
    .A(_01544_),
    .B(_05583_),
    .Y(_05584_)
  );
  NAND _13876_ (
    .A(_01521_),
    .B(_05582_),
    .Y(_05585_)
  );
  NAND _13877_ (
    .A(_05584_),
    .B(_05585_),
    .Y(_05586_)
  );
  OR _13878_ (
    .A(\data_i[7] ),
    .B(_01544_),
    .Y(_05587_)
  );
  AND _13879_ (
    .A(MemWrite_i),
    .B(_05587_),
    .Y(_05588_)
  );
  NAND _13880_ (
    .A(_05586_),
    .B(_05588_),
    .Y(_05590_)
  );
  NAND _13881_ (
    .A(_05575_),
    .B(_05590_),
    .Y(_00047_)
  );
  NAND _13882_ (
    .A(\memory[13][0] ),
    .B(_05361_),
    .Y(_05591_)
  );
  OR _13883_ (
    .A(\memory[13][0] ),
    .B(_01578_),
    .Y(_05592_)
  );
  OR _13884_ (
    .A(\data_i[24] ),
    .B(_01579_),
    .Y(_05593_)
  );
  NAND _13885_ (
    .A(_05592_),
    .B(_05593_),
    .Y(_05594_)
  );
  NAND _13886_ (
    .A(_01576_),
    .B(_05594_),
    .Y(_05595_)
  );
  OR _13887_ (
    .A(\data_i[16] ),
    .B(_01576_),
    .Y(_05596_)
  );
  AND _13888_ (
    .A(_05595_),
    .B(_05596_),
    .Y(_05597_)
  );
  NAND _13889_ (
    .A(\data_i[8] ),
    .B(_01458_),
    .Y(_05598_)
  );
  AND _13890_ (
    .A(_01521_),
    .B(_05598_),
    .Y(_05600_)
  );
  NAND _13891_ (
    .A(_01459_),
    .B(_05597_),
    .Y(_05601_)
  );
  NAND _13892_ (
    .A(_05600_),
    .B(_05601_),
    .Y(_05602_)
  );
  OR _13893_ (
    .A(\data_i[0] ),
    .B(_01521_),
    .Y(_05603_)
  );
  AND _13894_ (
    .A(MemWrite_i),
    .B(_05603_),
    .Y(_05604_)
  );
  NAND _13895_ (
    .A(_05602_),
    .B(_05604_),
    .Y(_05605_)
  );
  NAND _13896_ (
    .A(_05591_),
    .B(_05605_),
    .Y(_00032_)
  );
  NAND _13897_ (
    .A(\memory[13][1] ),
    .B(_05361_),
    .Y(_05606_)
  );
  OR _13898_ (
    .A(\memory[13][1] ),
    .B(_01578_),
    .Y(_05607_)
  );
  OR _13899_ (
    .A(\data_i[25] ),
    .B(_01579_),
    .Y(_05608_)
  );
  NAND _13900_ (
    .A(_05607_),
    .B(_05608_),
    .Y(_05610_)
  );
  NAND _13901_ (
    .A(_01576_),
    .B(_05610_),
    .Y(_05611_)
  );
  OR _13902_ (
    .A(\data_i[17] ),
    .B(_01576_),
    .Y(_05612_)
  );
  AND _13903_ (
    .A(_05611_),
    .B(_05612_),
    .Y(_05613_)
  );
  NAND _13904_ (
    .A(\data_i[9] ),
    .B(_01458_),
    .Y(_05614_)
  );
  AND _13905_ (
    .A(_01521_),
    .B(_05614_),
    .Y(_05615_)
  );
  NAND _13906_ (
    .A(_01459_),
    .B(_05613_),
    .Y(_05616_)
  );
  NAND _13907_ (
    .A(_05615_),
    .B(_05616_),
    .Y(_05617_)
  );
  OR _13908_ (
    .A(\data_i[1] ),
    .B(_01521_),
    .Y(_05618_)
  );
  AND _13909_ (
    .A(MemWrite_i),
    .B(_05618_),
    .Y(_05619_)
  );
  NAND _13910_ (
    .A(_05617_),
    .B(_05619_),
    .Y(_05621_)
  );
  NAND _13911_ (
    .A(_05606_),
    .B(_05621_),
    .Y(_00033_)
  );
  NAND _13912_ (
    .A(\memory[13][2] ),
    .B(_05361_),
    .Y(_05622_)
  );
  OR _13913_ (
    .A(\memory[13][2] ),
    .B(_01578_),
    .Y(_05623_)
  );
  OR _13914_ (
    .A(\data_i[26] ),
    .B(_01579_),
    .Y(_05624_)
  );
  NAND _13915_ (
    .A(_05623_),
    .B(_05624_),
    .Y(_05625_)
  );
  NAND _13916_ (
    .A(_01576_),
    .B(_05625_),
    .Y(_05626_)
  );
  OR _13917_ (
    .A(\data_i[18] ),
    .B(_01576_),
    .Y(_05627_)
  );
  AND _13918_ (
    .A(_05626_),
    .B(_05627_),
    .Y(_05628_)
  );
  NAND _13919_ (
    .A(\data_i[10] ),
    .B(_01458_),
    .Y(_05629_)
  );
  AND _13920_ (
    .A(_01521_),
    .B(_05629_),
    .Y(_05631_)
  );
  NAND _13921_ (
    .A(_01459_),
    .B(_05628_),
    .Y(_05632_)
  );
  NAND _13922_ (
    .A(_05631_),
    .B(_05632_),
    .Y(_05633_)
  );
  OR _13923_ (
    .A(\data_i[2] ),
    .B(_01521_),
    .Y(_05634_)
  );
  AND _13924_ (
    .A(MemWrite_i),
    .B(_05634_),
    .Y(_05635_)
  );
  NAND _13925_ (
    .A(_05633_),
    .B(_05635_),
    .Y(_05636_)
  );
  NAND _13926_ (
    .A(_05622_),
    .B(_05636_),
    .Y(_00034_)
  );
  NAND _13927_ (
    .A(\memory[13][3] ),
    .B(_05361_),
    .Y(_05637_)
  );
  OR _13928_ (
    .A(\memory[13][3] ),
    .B(_01578_),
    .Y(_05638_)
  );
  OR _13929_ (
    .A(\data_i[27] ),
    .B(_01579_),
    .Y(_05639_)
  );
  NAND _13930_ (
    .A(_05638_),
    .B(_05639_),
    .Y(_05641_)
  );
  NAND _13931_ (
    .A(_01576_),
    .B(_05641_),
    .Y(_05642_)
  );
  OR _13932_ (
    .A(\data_i[19] ),
    .B(_01576_),
    .Y(_05643_)
  );
  AND _13933_ (
    .A(_05642_),
    .B(_05643_),
    .Y(_05644_)
  );
  NAND _13934_ (
    .A(\data_i[11] ),
    .B(_01458_),
    .Y(_05645_)
  );
  AND _13935_ (
    .A(_01521_),
    .B(_05645_),
    .Y(_05646_)
  );
  NAND _13936_ (
    .A(_01459_),
    .B(_05644_),
    .Y(_05647_)
  );
  NAND _13937_ (
    .A(_05646_),
    .B(_05647_),
    .Y(_05648_)
  );
  OR _13938_ (
    .A(\data_i[3] ),
    .B(_01521_),
    .Y(_05649_)
  );
  AND _13939_ (
    .A(MemWrite_i),
    .B(_05649_),
    .Y(_05650_)
  );
  NAND _13940_ (
    .A(_05648_),
    .B(_05650_),
    .Y(_05652_)
  );
  NAND _13941_ (
    .A(_05637_),
    .B(_05652_),
    .Y(_00035_)
  );
  NAND _13942_ (
    .A(\memory[13][4] ),
    .B(_05361_),
    .Y(_05653_)
  );
  OR _13943_ (
    .A(\memory[13][4] ),
    .B(_01578_),
    .Y(_05654_)
  );
  OR _13944_ (
    .A(\data_i[28] ),
    .B(_01579_),
    .Y(_05655_)
  );
  NAND _13945_ (
    .A(_05654_),
    .B(_05655_),
    .Y(_05656_)
  );
  NAND _13946_ (
    .A(_01576_),
    .B(_05656_),
    .Y(_05657_)
  );
  OR _13947_ (
    .A(\data_i[20] ),
    .B(_01576_),
    .Y(_05658_)
  );
  AND _13948_ (
    .A(_05657_),
    .B(_05658_),
    .Y(_05659_)
  );
  NAND _13949_ (
    .A(\data_i[12] ),
    .B(_01458_),
    .Y(_05660_)
  );
  AND _13950_ (
    .A(_01521_),
    .B(_05660_),
    .Y(_05662_)
  );
  NAND _13951_ (
    .A(_01459_),
    .B(_05659_),
    .Y(_05663_)
  );
  NAND _13952_ (
    .A(_05662_),
    .B(_05663_),
    .Y(_05664_)
  );
  OR _13953_ (
    .A(\data_i[4] ),
    .B(_01521_),
    .Y(_05665_)
  );
  AND _13954_ (
    .A(MemWrite_i),
    .B(_05665_),
    .Y(_05666_)
  );
  NAND _13955_ (
    .A(_05664_),
    .B(_05666_),
    .Y(_05667_)
  );
  NAND _13956_ (
    .A(_05653_),
    .B(_05667_),
    .Y(_00036_)
  );
  NAND _13957_ (
    .A(\memory[13][5] ),
    .B(_05361_),
    .Y(_05668_)
  );
  OR _13958_ (
    .A(\memory[13][5] ),
    .B(_01578_),
    .Y(_05669_)
  );
  OR _13959_ (
    .A(\data_i[29] ),
    .B(_01579_),
    .Y(_05670_)
  );
  NAND _13960_ (
    .A(_05669_),
    .B(_05670_),
    .Y(_05672_)
  );
  NAND _13961_ (
    .A(_01576_),
    .B(_05672_),
    .Y(_05673_)
  );
  OR _13962_ (
    .A(\data_i[21] ),
    .B(_01576_),
    .Y(_05674_)
  );
  AND _13963_ (
    .A(_05673_),
    .B(_05674_),
    .Y(_05675_)
  );
  NAND _13964_ (
    .A(\data_i[13] ),
    .B(_01458_),
    .Y(_05676_)
  );
  AND _13965_ (
    .A(_01521_),
    .B(_05676_),
    .Y(_05677_)
  );
  NAND _13966_ (
    .A(_01459_),
    .B(_05675_),
    .Y(_05678_)
  );
  NAND _13967_ (
    .A(_05677_),
    .B(_05678_),
    .Y(_05679_)
  );
  OR _13968_ (
    .A(\data_i[5] ),
    .B(_01521_),
    .Y(_05680_)
  );
  AND _13969_ (
    .A(MemWrite_i),
    .B(_05680_),
    .Y(_05681_)
  );
  NAND _13970_ (
    .A(_05679_),
    .B(_05681_),
    .Y(_05683_)
  );
  NAND _13971_ (
    .A(_05668_),
    .B(_05683_),
    .Y(_00037_)
  );
  NAND _13972_ (
    .A(\memory[13][6] ),
    .B(_05361_),
    .Y(_05684_)
  );
  OR _13973_ (
    .A(\memory[13][6] ),
    .B(_01578_),
    .Y(_05685_)
  );
  OR _13974_ (
    .A(\data_i[30] ),
    .B(_01579_),
    .Y(_05686_)
  );
  NAND _13975_ (
    .A(_05685_),
    .B(_05686_),
    .Y(_05687_)
  );
  NAND _13976_ (
    .A(_01576_),
    .B(_05687_),
    .Y(_05688_)
  );
  OR _13977_ (
    .A(\data_i[22] ),
    .B(_01576_),
    .Y(_05689_)
  );
  AND _13978_ (
    .A(_05688_),
    .B(_05689_),
    .Y(_05690_)
  );
  NAND _13979_ (
    .A(\data_i[14] ),
    .B(_01458_),
    .Y(_05691_)
  );
  AND _13980_ (
    .A(_01521_),
    .B(_05691_),
    .Y(_05693_)
  );
  NAND _13981_ (
    .A(_01459_),
    .B(_05690_),
    .Y(_05694_)
  );
  NAND _13982_ (
    .A(_05693_),
    .B(_05694_),
    .Y(_05695_)
  );
  OR _13983_ (
    .A(\data_i[6] ),
    .B(_01521_),
    .Y(_05696_)
  );
  AND _13984_ (
    .A(MemWrite_i),
    .B(_05696_),
    .Y(_05697_)
  );
  NAND _13985_ (
    .A(_05695_),
    .B(_05697_),
    .Y(_05698_)
  );
  NAND _13986_ (
    .A(_05684_),
    .B(_05698_),
    .Y(_00038_)
  );
  NAND _13987_ (
    .A(\memory[13][7] ),
    .B(_05361_),
    .Y(_05699_)
  );
  OR _13988_ (
    .A(\memory[13][7] ),
    .B(_01578_),
    .Y(_05700_)
  );
  OR _13989_ (
    .A(\data_i[31] ),
    .B(_01579_),
    .Y(_05701_)
  );
  NAND _13990_ (
    .A(_05700_),
    .B(_05701_),
    .Y(_05703_)
  );
  NAND _13991_ (
    .A(_01576_),
    .B(_05703_),
    .Y(_05704_)
  );
  OR _13992_ (
    .A(\data_i[23] ),
    .B(_01576_),
    .Y(_05705_)
  );
  AND _13993_ (
    .A(_05704_),
    .B(_05705_),
    .Y(_05706_)
  );
  NAND _13994_ (
    .A(\data_i[15] ),
    .B(_01458_),
    .Y(_05707_)
  );
  AND _13995_ (
    .A(_01521_),
    .B(_05707_),
    .Y(_05708_)
  );
  NAND _13996_ (
    .A(_01459_),
    .B(_05706_),
    .Y(_05709_)
  );
  NAND _13997_ (
    .A(_05708_),
    .B(_05709_),
    .Y(_05710_)
  );
  OR _13998_ (
    .A(\data_i[7] ),
    .B(_01521_),
    .Y(_05711_)
  );
  AND _13999_ (
    .A(MemWrite_i),
    .B(_05711_),
    .Y(_05712_)
  );
  NAND _14000_ (
    .A(_05710_),
    .B(_05712_),
    .Y(_05714_)
  );
  NAND _14001_ (
    .A(_05699_),
    .B(_05714_),
    .Y(_00039_)
  );
  NAND _14002_ (
    .A(\memory[12][0] ),
    .B(_05361_),
    .Y(_05715_)
  );
  OR _14003_ (
    .A(\memory[12][0] ),
    .B(_01495_),
    .Y(_05716_)
  );
  OR _14004_ (
    .A(\data_i[24] ),
    .B(_01496_),
    .Y(_05717_)
  );
  NAND _14005_ (
    .A(_05716_),
    .B(_05717_),
    .Y(_05718_)
  );
  NAND _14006_ (
    .A(_01579_),
    .B(_05718_),
    .Y(_05719_)
  );
  OR _14007_ (
    .A(\data_i[16] ),
    .B(_01579_),
    .Y(_05720_)
  );
  AND _14008_ (
    .A(_05719_),
    .B(_05720_),
    .Y(_05721_)
  );
  NAND _14009_ (
    .A(\data_i[8] ),
    .B(_01575_),
    .Y(_05722_)
  );
  AND _14010_ (
    .A(_01459_),
    .B(_05722_),
    .Y(_05724_)
  );
  NAND _14011_ (
    .A(_01576_),
    .B(_05721_),
    .Y(_05725_)
  );
  NAND _14012_ (
    .A(_05724_),
    .B(_05725_),
    .Y(_05726_)
  );
  OR _14013_ (
    .A(\data_i[0] ),
    .B(_01459_),
    .Y(_05727_)
  );
  AND _14014_ (
    .A(MemWrite_i),
    .B(_05727_),
    .Y(_05728_)
  );
  NAND _14015_ (
    .A(_05726_),
    .B(_05728_),
    .Y(_05729_)
  );
  NAND _14016_ (
    .A(_05715_),
    .B(_05729_),
    .Y(_00024_)
  );
  NAND _14017_ (
    .A(\memory[12][1] ),
    .B(_05361_),
    .Y(_05730_)
  );
  OR _14018_ (
    .A(\memory[12][1] ),
    .B(_01495_),
    .Y(_05731_)
  );
  OR _14019_ (
    .A(\data_i[25] ),
    .B(_01496_),
    .Y(_05732_)
  );
  NAND _14020_ (
    .A(_05731_),
    .B(_05732_),
    .Y(_05734_)
  );
  NAND _14021_ (
    .A(_01579_),
    .B(_05734_),
    .Y(_05735_)
  );
  OR _14022_ (
    .A(\data_i[17] ),
    .B(_01579_),
    .Y(_05736_)
  );
  AND _14023_ (
    .A(_05735_),
    .B(_05736_),
    .Y(_05737_)
  );
  NAND _14024_ (
    .A(\data_i[9] ),
    .B(_01575_),
    .Y(_05738_)
  );
  AND _14025_ (
    .A(_01459_),
    .B(_05738_),
    .Y(_05739_)
  );
  NAND _14026_ (
    .A(_01576_),
    .B(_05737_),
    .Y(_05740_)
  );
  NAND _14027_ (
    .A(_05739_),
    .B(_05740_),
    .Y(_05741_)
  );
  OR _14028_ (
    .A(\data_i[1] ),
    .B(_01459_),
    .Y(_05742_)
  );
  AND _14029_ (
    .A(MemWrite_i),
    .B(_05742_),
    .Y(_05743_)
  );
  NAND _14030_ (
    .A(_05741_),
    .B(_05743_),
    .Y(_05745_)
  );
  NAND _14031_ (
    .A(_05730_),
    .B(_05745_),
    .Y(_00025_)
  );
  NAND _14032_ (
    .A(\memory[12][2] ),
    .B(_05361_),
    .Y(_05746_)
  );
  OR _14033_ (
    .A(\memory[12][2] ),
    .B(_01495_),
    .Y(_05747_)
  );
  OR _14034_ (
    .A(\data_i[26] ),
    .B(_01496_),
    .Y(_05748_)
  );
  NAND _14035_ (
    .A(_05747_),
    .B(_05748_),
    .Y(_05749_)
  );
  NAND _14036_ (
    .A(_01579_),
    .B(_05749_),
    .Y(_05750_)
  );
  OR _14037_ (
    .A(\data_i[18] ),
    .B(_01579_),
    .Y(_05751_)
  );
  AND _14038_ (
    .A(_05750_),
    .B(_05751_),
    .Y(_05752_)
  );
  NAND _14039_ (
    .A(\data_i[10] ),
    .B(_01575_),
    .Y(_05753_)
  );
  AND _14040_ (
    .A(_01459_),
    .B(_05753_),
    .Y(_05755_)
  );
  NAND _14041_ (
    .A(_01576_),
    .B(_05752_),
    .Y(_05756_)
  );
  NAND _14042_ (
    .A(_05755_),
    .B(_05756_),
    .Y(_05757_)
  );
  OR _14043_ (
    .A(\data_i[2] ),
    .B(_01459_),
    .Y(_05758_)
  );
  AND _14044_ (
    .A(MemWrite_i),
    .B(_05758_),
    .Y(_05759_)
  );
  NAND _14045_ (
    .A(_05757_),
    .B(_05759_),
    .Y(_05760_)
  );
  NAND _14046_ (
    .A(_05746_),
    .B(_05760_),
    .Y(_00026_)
  );
  NAND _14047_ (
    .A(\memory[12][3] ),
    .B(_05361_),
    .Y(_05761_)
  );
  OR _14048_ (
    .A(\memory[12][3] ),
    .B(_01495_),
    .Y(_05762_)
  );
  OR _14049_ (
    .A(\data_i[27] ),
    .B(_01496_),
    .Y(_05763_)
  );
  NAND _14050_ (
    .A(_05762_),
    .B(_05763_),
    .Y(_05765_)
  );
  NAND _14051_ (
    .A(_01579_),
    .B(_05765_),
    .Y(_05766_)
  );
  OR _14052_ (
    .A(\data_i[19] ),
    .B(_01579_),
    .Y(_05767_)
  );
  AND _14053_ (
    .A(_05766_),
    .B(_05767_),
    .Y(_05768_)
  );
  NAND _14054_ (
    .A(\data_i[11] ),
    .B(_01575_),
    .Y(_05769_)
  );
  AND _14055_ (
    .A(_01459_),
    .B(_05769_),
    .Y(_05770_)
  );
  NAND _14056_ (
    .A(_01576_),
    .B(_05768_),
    .Y(_05771_)
  );
  NAND _14057_ (
    .A(_05770_),
    .B(_05771_),
    .Y(_05772_)
  );
  OR _14058_ (
    .A(\data_i[3] ),
    .B(_01459_),
    .Y(_05773_)
  );
  AND _14059_ (
    .A(MemWrite_i),
    .B(_05773_),
    .Y(_05774_)
  );
  NAND _14060_ (
    .A(_05772_),
    .B(_05774_),
    .Y(_05776_)
  );
  NAND _14061_ (
    .A(_05761_),
    .B(_05776_),
    .Y(_00027_)
  );
  NAND _14062_ (
    .A(\memory[12][4] ),
    .B(_05361_),
    .Y(_05777_)
  );
  OR _14063_ (
    .A(\memory[12][4] ),
    .B(_01495_),
    .Y(_05778_)
  );
  OR _14064_ (
    .A(\data_i[28] ),
    .B(_01496_),
    .Y(_05779_)
  );
  NAND _14065_ (
    .A(_05778_),
    .B(_05779_),
    .Y(_05780_)
  );
  NAND _14066_ (
    .A(_01579_),
    .B(_05780_),
    .Y(_05781_)
  );
  OR _14067_ (
    .A(\data_i[20] ),
    .B(_01579_),
    .Y(_05782_)
  );
  AND _14068_ (
    .A(_05781_),
    .B(_05782_),
    .Y(_05783_)
  );
  NAND _14069_ (
    .A(\data_i[12] ),
    .B(_01575_),
    .Y(_05784_)
  );
  AND _14070_ (
    .A(_01459_),
    .B(_05784_),
    .Y(_05786_)
  );
  NAND _14071_ (
    .A(_01576_),
    .B(_05783_),
    .Y(_05787_)
  );
  NAND _14072_ (
    .A(_05786_),
    .B(_05787_),
    .Y(_05788_)
  );
  OR _14073_ (
    .A(\data_i[4] ),
    .B(_01459_),
    .Y(_05789_)
  );
  AND _14074_ (
    .A(MemWrite_i),
    .B(_05789_),
    .Y(_05790_)
  );
  NAND _14075_ (
    .A(_05788_),
    .B(_05790_),
    .Y(_05791_)
  );
  NAND _14076_ (
    .A(_05777_),
    .B(_05791_),
    .Y(_00028_)
  );
  NAND _14077_ (
    .A(\memory[12][5] ),
    .B(_05361_),
    .Y(_05792_)
  );
  OR _14078_ (
    .A(\memory[12][5] ),
    .B(_01495_),
    .Y(_05793_)
  );
  OR _14079_ (
    .A(\data_i[29] ),
    .B(_01496_),
    .Y(_05794_)
  );
  NAND _14080_ (
    .A(_05793_),
    .B(_05794_),
    .Y(_05796_)
  );
  NAND _14081_ (
    .A(_01579_),
    .B(_05796_),
    .Y(_05797_)
  );
  OR _14082_ (
    .A(\data_i[21] ),
    .B(_01579_),
    .Y(_05798_)
  );
  AND _14083_ (
    .A(_05797_),
    .B(_05798_),
    .Y(_05799_)
  );
  NAND _14084_ (
    .A(\data_i[13] ),
    .B(_01575_),
    .Y(_05800_)
  );
  AND _14085_ (
    .A(_01459_),
    .B(_05800_),
    .Y(_05801_)
  );
  NAND _14086_ (
    .A(_01576_),
    .B(_05799_),
    .Y(_05802_)
  );
  NAND _14087_ (
    .A(_05801_),
    .B(_05802_),
    .Y(_05803_)
  );
  OR _14088_ (
    .A(\data_i[5] ),
    .B(_01459_),
    .Y(_05804_)
  );
  AND _14089_ (
    .A(MemWrite_i),
    .B(_05804_),
    .Y(_05805_)
  );
  NAND _14090_ (
    .A(_05803_),
    .B(_05805_),
    .Y(_05807_)
  );
  NAND _14091_ (
    .A(_05792_),
    .B(_05807_),
    .Y(_00029_)
  );
  NAND _14092_ (
    .A(\memory[12][6] ),
    .B(_05361_),
    .Y(_05808_)
  );
  OR _14093_ (
    .A(\memory[12][6] ),
    .B(_01495_),
    .Y(_05809_)
  );
  OR _14094_ (
    .A(\data_i[30] ),
    .B(_01496_),
    .Y(_05810_)
  );
  NAND _14095_ (
    .A(_05809_),
    .B(_05810_),
    .Y(_05811_)
  );
  NAND _14096_ (
    .A(_01579_),
    .B(_05811_),
    .Y(_05812_)
  );
  OR _14097_ (
    .A(\data_i[22] ),
    .B(_01579_),
    .Y(_05813_)
  );
  AND _14098_ (
    .A(_05812_),
    .B(_05813_),
    .Y(_05814_)
  );
  NAND _14099_ (
    .A(\data_i[14] ),
    .B(_01575_),
    .Y(_05815_)
  );
  AND _14100_ (
    .A(_01459_),
    .B(_05815_),
    .Y(_05817_)
  );
  NAND _14101_ (
    .A(_01576_),
    .B(_05814_),
    .Y(_05818_)
  );
  NAND _14102_ (
    .A(_05817_),
    .B(_05818_),
    .Y(_05819_)
  );
  OR _14103_ (
    .A(\data_i[6] ),
    .B(_01459_),
    .Y(_05820_)
  );
  AND _14104_ (
    .A(MemWrite_i),
    .B(_05820_),
    .Y(_05821_)
  );
  NAND _14105_ (
    .A(_05819_),
    .B(_05821_),
    .Y(_05822_)
  );
  NAND _14106_ (
    .A(_05808_),
    .B(_05822_),
    .Y(_00030_)
  );
  NAND _14107_ (
    .A(\memory[12][7] ),
    .B(_05361_),
    .Y(_05823_)
  );
  OR _14108_ (
    .A(\memory[12][7] ),
    .B(_01495_),
    .Y(_05824_)
  );
  OR _14109_ (
    .A(\data_i[31] ),
    .B(_01496_),
    .Y(_05825_)
  );
  NAND _14110_ (
    .A(_05824_),
    .B(_05825_),
    .Y(_05827_)
  );
  NAND _14111_ (
    .A(_01579_),
    .B(_05827_),
    .Y(_05828_)
  );
  OR _14112_ (
    .A(\data_i[23] ),
    .B(_01579_),
    .Y(_05829_)
  );
  AND _14113_ (
    .A(_05828_),
    .B(_05829_),
    .Y(_05830_)
  );
  NAND _14114_ (
    .A(\data_i[15] ),
    .B(_01575_),
    .Y(_05831_)
  );
  AND _14115_ (
    .A(_01459_),
    .B(_05831_),
    .Y(_05832_)
  );
  NAND _14116_ (
    .A(_01576_),
    .B(_05830_),
    .Y(_05833_)
  );
  NAND _14117_ (
    .A(_05832_),
    .B(_05833_),
    .Y(_05834_)
  );
  OR _14118_ (
    .A(\data_i[7] ),
    .B(_01459_),
    .Y(_05835_)
  );
  AND _14119_ (
    .A(MemWrite_i),
    .B(_05835_),
    .Y(_05836_)
  );
  NAND _14120_ (
    .A(_05834_),
    .B(_05836_),
    .Y(_05838_)
  );
  NAND _14121_ (
    .A(_05823_),
    .B(_05838_),
    .Y(_00031_)
  );
  NAND _14122_ (
    .A(\memory[11][0] ),
    .B(_05361_),
    .Y(_05839_)
  );
  OR _14123_ (
    .A(\memory[11][0] ),
    .B(_01527_),
    .Y(_05840_)
  );
  OR _14124_ (
    .A(\data_i[24] ),
    .B(_01528_),
    .Y(_05841_)
  );
  NAND _14125_ (
    .A(_05840_),
    .B(_05841_),
    .Y(_05842_)
  );
  NAND _14126_ (
    .A(_01496_),
    .B(_05842_),
    .Y(_05843_)
  );
  OR _14127_ (
    .A(\data_i[16] ),
    .B(_01496_),
    .Y(_05844_)
  );
  AND _14128_ (
    .A(_05843_),
    .B(_05844_),
    .Y(_05845_)
  );
  NAND _14129_ (
    .A(\data_i[8] ),
    .B(_01578_),
    .Y(_05846_)
  );
  AND _14130_ (
    .A(_01576_),
    .B(_05846_),
    .Y(_05848_)
  );
  NAND _14131_ (
    .A(_01579_),
    .B(_05845_),
    .Y(_05849_)
  );
  NAND _14132_ (
    .A(_05848_),
    .B(_05849_),
    .Y(_05850_)
  );
  OR _14133_ (
    .A(\data_i[0] ),
    .B(_01576_),
    .Y(_05851_)
  );
  AND _14134_ (
    .A(MemWrite_i),
    .B(_05851_),
    .Y(_05852_)
  );
  NAND _14135_ (
    .A(_05850_),
    .B(_05852_),
    .Y(_05853_)
  );
  NAND _14136_ (
    .A(_05839_),
    .B(_05853_),
    .Y(_00016_)
  );
  NAND _14137_ (
    .A(\memory[11][1] ),
    .B(_05361_),
    .Y(_05854_)
  );
  OR _14138_ (
    .A(\memory[11][1] ),
    .B(_01527_),
    .Y(_05855_)
  );
  OR _14139_ (
    .A(\data_i[25] ),
    .B(_01528_),
    .Y(_05856_)
  );
  NAND _14140_ (
    .A(_05855_),
    .B(_05856_),
    .Y(_05858_)
  );
  NAND _14141_ (
    .A(_01496_),
    .B(_05858_),
    .Y(_05859_)
  );
  OR _14142_ (
    .A(\data_i[17] ),
    .B(_01496_),
    .Y(_05860_)
  );
  AND _14143_ (
    .A(_05859_),
    .B(_05860_),
    .Y(_05861_)
  );
  NAND _14144_ (
    .A(\data_i[9] ),
    .B(_01578_),
    .Y(_05862_)
  );
  AND _14145_ (
    .A(_01576_),
    .B(_05862_),
    .Y(_05863_)
  );
  NAND _14146_ (
    .A(_01579_),
    .B(_05861_),
    .Y(_05864_)
  );
  NAND _14147_ (
    .A(_05863_),
    .B(_05864_),
    .Y(_05865_)
  );
  OR _14148_ (
    .A(\data_i[1] ),
    .B(_01576_),
    .Y(_05866_)
  );
  AND _14149_ (
    .A(MemWrite_i),
    .B(_05866_),
    .Y(_05867_)
  );
  NAND _14150_ (
    .A(_05865_),
    .B(_05867_),
    .Y(_05869_)
  );
  NAND _14151_ (
    .A(_05854_),
    .B(_05869_),
    .Y(_00017_)
  );
  NAND _14152_ (
    .A(\memory[11][2] ),
    .B(_05361_),
    .Y(_05870_)
  );
  OR _14153_ (
    .A(\memory[11][2] ),
    .B(_01527_),
    .Y(_05871_)
  );
  OR _14154_ (
    .A(\data_i[26] ),
    .B(_01528_),
    .Y(_05872_)
  );
  NAND _14155_ (
    .A(_05871_),
    .B(_05872_),
    .Y(_05873_)
  );
  NAND _14156_ (
    .A(_01496_),
    .B(_05873_),
    .Y(_05874_)
  );
  OR _14157_ (
    .A(\data_i[18] ),
    .B(_01496_),
    .Y(_05875_)
  );
  AND _14158_ (
    .A(_05874_),
    .B(_05875_),
    .Y(_05876_)
  );
  NAND _14159_ (
    .A(\data_i[10] ),
    .B(_01578_),
    .Y(_05877_)
  );
  AND _14160_ (
    .A(_01576_),
    .B(_05877_),
    .Y(_05879_)
  );
  NAND _14161_ (
    .A(_01579_),
    .B(_05876_),
    .Y(_05880_)
  );
  NAND _14162_ (
    .A(_05879_),
    .B(_05880_),
    .Y(_05881_)
  );
  OR _14163_ (
    .A(\data_i[2] ),
    .B(_01576_),
    .Y(_05882_)
  );
  AND _14164_ (
    .A(MemWrite_i),
    .B(_05882_),
    .Y(_05883_)
  );
  NAND _14165_ (
    .A(_05881_),
    .B(_05883_),
    .Y(_05884_)
  );
  NAND _14166_ (
    .A(_05870_),
    .B(_05884_),
    .Y(_00018_)
  );
  NAND _14167_ (
    .A(\memory[11][3] ),
    .B(_05361_),
    .Y(_05885_)
  );
  OR _14168_ (
    .A(\memory[11][3] ),
    .B(_01527_),
    .Y(_05886_)
  );
  OR _14169_ (
    .A(\data_i[27] ),
    .B(_01528_),
    .Y(_05887_)
  );
  NAND _14170_ (
    .A(_05886_),
    .B(_05887_),
    .Y(_05889_)
  );
  NAND _14171_ (
    .A(_01496_),
    .B(_05889_),
    .Y(_05890_)
  );
  OR _14172_ (
    .A(\data_i[19] ),
    .B(_01496_),
    .Y(_05891_)
  );
  AND _14173_ (
    .A(_05890_),
    .B(_05891_),
    .Y(_05892_)
  );
  NAND _14174_ (
    .A(\data_i[11] ),
    .B(_01578_),
    .Y(_05893_)
  );
  AND _14175_ (
    .A(_01576_),
    .B(_05893_),
    .Y(_05894_)
  );
  NAND _14176_ (
    .A(_01579_),
    .B(_05892_),
    .Y(_05895_)
  );
  NAND _14177_ (
    .A(_05894_),
    .B(_05895_),
    .Y(_05896_)
  );
  OR _14178_ (
    .A(\data_i[3] ),
    .B(_01576_),
    .Y(_05897_)
  );
  AND _14179_ (
    .A(MemWrite_i),
    .B(_05897_),
    .Y(_05898_)
  );
  NAND _14180_ (
    .A(_05896_),
    .B(_05898_),
    .Y(_05900_)
  );
  NAND _14181_ (
    .A(_05885_),
    .B(_05900_),
    .Y(_00019_)
  );
  NAND _14182_ (
    .A(\memory[11][4] ),
    .B(_05361_),
    .Y(_05901_)
  );
  OR _14183_ (
    .A(\memory[11][4] ),
    .B(_01527_),
    .Y(_05902_)
  );
  OR _14184_ (
    .A(\data_i[28] ),
    .B(_01528_),
    .Y(_05903_)
  );
  NAND _14185_ (
    .A(_05902_),
    .B(_05903_),
    .Y(_05904_)
  );
  NAND _14186_ (
    .A(_01496_),
    .B(_05904_),
    .Y(_05905_)
  );
  OR _14187_ (
    .A(\data_i[20] ),
    .B(_01496_),
    .Y(_05906_)
  );
  AND _14188_ (
    .A(_05905_),
    .B(_05906_),
    .Y(_05907_)
  );
  NAND _14189_ (
    .A(\data_i[12] ),
    .B(_01578_),
    .Y(_05908_)
  );
  AND _14190_ (
    .A(_01576_),
    .B(_05908_),
    .Y(_05910_)
  );
  NAND _14191_ (
    .A(_01579_),
    .B(_05907_),
    .Y(_05911_)
  );
  NAND _14192_ (
    .A(_05910_),
    .B(_05911_),
    .Y(_05912_)
  );
  OR _14193_ (
    .A(\data_i[4] ),
    .B(_01576_),
    .Y(_05913_)
  );
  AND _14194_ (
    .A(MemWrite_i),
    .B(_05913_),
    .Y(_05914_)
  );
  NAND _14195_ (
    .A(_05912_),
    .B(_05914_),
    .Y(_05915_)
  );
  NAND _14196_ (
    .A(_05901_),
    .B(_05915_),
    .Y(_00020_)
  );
  NAND _14197_ (
    .A(\memory[11][5] ),
    .B(_05361_),
    .Y(_05916_)
  );
  OR _14198_ (
    .A(\memory[11][5] ),
    .B(_01527_),
    .Y(_05917_)
  );
  OR _14199_ (
    .A(\data_i[29] ),
    .B(_01528_),
    .Y(_05918_)
  );
  NAND _14200_ (
    .A(_05917_),
    .B(_05918_),
    .Y(_05920_)
  );
  NAND _14201_ (
    .A(_01496_),
    .B(_05920_),
    .Y(_05921_)
  );
  OR _14202_ (
    .A(\data_i[21] ),
    .B(_01496_),
    .Y(_05922_)
  );
  AND _14203_ (
    .A(_05921_),
    .B(_05922_),
    .Y(_05923_)
  );
  NAND _14204_ (
    .A(\data_i[13] ),
    .B(_01578_),
    .Y(_05924_)
  );
  AND _14205_ (
    .A(_01576_),
    .B(_05924_),
    .Y(_05925_)
  );
  NAND _14206_ (
    .A(_01579_),
    .B(_05923_),
    .Y(_05926_)
  );
  NAND _14207_ (
    .A(_05925_),
    .B(_05926_),
    .Y(_05927_)
  );
  OR _14208_ (
    .A(\data_i[5] ),
    .B(_01576_),
    .Y(_05928_)
  );
  AND _14209_ (
    .A(MemWrite_i),
    .B(_05928_),
    .Y(_05929_)
  );
  NAND _14210_ (
    .A(_05927_),
    .B(_05929_),
    .Y(_05931_)
  );
  NAND _14211_ (
    .A(_05916_),
    .B(_05931_),
    .Y(_00021_)
  );
  NAND _14212_ (
    .A(\memory[11][6] ),
    .B(_05361_),
    .Y(_05932_)
  );
  OR _14213_ (
    .A(\memory[11][6] ),
    .B(_01527_),
    .Y(_05933_)
  );
  OR _14214_ (
    .A(\data_i[30] ),
    .B(_01528_),
    .Y(_05934_)
  );
  NAND _14215_ (
    .A(_05933_),
    .B(_05934_),
    .Y(_05935_)
  );
  NAND _14216_ (
    .A(_01496_),
    .B(_05935_),
    .Y(_05936_)
  );
  OR _14217_ (
    .A(\data_i[22] ),
    .B(_01496_),
    .Y(_05937_)
  );
  AND _14218_ (
    .A(_05936_),
    .B(_05937_),
    .Y(_05938_)
  );
  NAND _14219_ (
    .A(\data_i[14] ),
    .B(_01578_),
    .Y(_05939_)
  );
  AND _14220_ (
    .A(_01576_),
    .B(_05939_),
    .Y(_05941_)
  );
  NAND _14221_ (
    .A(_01579_),
    .B(_05938_),
    .Y(_05942_)
  );
  NAND _14222_ (
    .A(_05941_),
    .B(_05942_),
    .Y(_05943_)
  );
  OR _14223_ (
    .A(\data_i[6] ),
    .B(_01576_),
    .Y(_05944_)
  );
  AND _14224_ (
    .A(MemWrite_i),
    .B(_05944_),
    .Y(_05945_)
  );
  NAND _14225_ (
    .A(_05943_),
    .B(_05945_),
    .Y(_05946_)
  );
  NAND _14226_ (
    .A(_05932_),
    .B(_05946_),
    .Y(_00022_)
  );
  NAND _14227_ (
    .A(\memory[11][7] ),
    .B(_05361_),
    .Y(_05947_)
  );
  OR _14228_ (
    .A(\memory[11][7] ),
    .B(_01527_),
    .Y(_05948_)
  );
  OR _14229_ (
    .A(\data_i[31] ),
    .B(_01528_),
    .Y(_05949_)
  );
  NAND _14230_ (
    .A(_05948_),
    .B(_05949_),
    .Y(_05951_)
  );
  NAND _14231_ (
    .A(_01496_),
    .B(_05951_),
    .Y(_05952_)
  );
  OR _14232_ (
    .A(\data_i[23] ),
    .B(_01496_),
    .Y(_05953_)
  );
  AND _14233_ (
    .A(_05952_),
    .B(_05953_),
    .Y(_05954_)
  );
  NAND _14234_ (
    .A(\data_i[15] ),
    .B(_01578_),
    .Y(_05955_)
  );
  AND _14235_ (
    .A(_01576_),
    .B(_05955_),
    .Y(_05956_)
  );
  NAND _14236_ (
    .A(_01579_),
    .B(_05954_),
    .Y(_05957_)
  );
  NAND _14237_ (
    .A(_05956_),
    .B(_05957_),
    .Y(_05958_)
  );
  OR _14238_ (
    .A(\data_i[7] ),
    .B(_01576_),
    .Y(_05959_)
  );
  AND _14239_ (
    .A(MemWrite_i),
    .B(_05959_),
    .Y(_05960_)
  );
  NAND _14240_ (
    .A(_05958_),
    .B(_05960_),
    .Y(_05962_)
  );
  NAND _14241_ (
    .A(_05947_),
    .B(_05962_),
    .Y(_00023_)
  );
  NAND _14242_ (
    .A(\memory[10][0] ),
    .B(_05361_),
    .Y(_05963_)
  );
  OR _14243_ (
    .A(\memory[10][0] ),
    .B(_01538_),
    .Y(_05964_)
  );
  OR _14244_ (
    .A(\data_i[24] ),
    .B(_01539_),
    .Y(_05965_)
  );
  NAND _14245_ (
    .A(_05964_),
    .B(_05965_),
    .Y(_05966_)
  );
  NAND _14246_ (
    .A(_01528_),
    .B(_05966_),
    .Y(_05967_)
  );
  OR _14247_ (
    .A(\data_i[16] ),
    .B(_01528_),
    .Y(_05968_)
  );
  AND _14248_ (
    .A(_05967_),
    .B(_05968_),
    .Y(_05969_)
  );
  NAND _14249_ (
    .A(\data_i[8] ),
    .B(_01495_),
    .Y(_05970_)
  );
  AND _14250_ (
    .A(_01579_),
    .B(_05970_),
    .Y(_05972_)
  );
  NAND _14251_ (
    .A(_01496_),
    .B(_05969_),
    .Y(_05973_)
  );
  NAND _14252_ (
    .A(_05972_),
    .B(_05973_),
    .Y(_05974_)
  );
  OR _14253_ (
    .A(\data_i[0] ),
    .B(_01579_),
    .Y(_05975_)
  );
  AND _14254_ (
    .A(MemWrite_i),
    .B(_05975_),
    .Y(_05976_)
  );
  NAND _14255_ (
    .A(_05974_),
    .B(_05976_),
    .Y(_05977_)
  );
  NAND _14256_ (
    .A(_05963_),
    .B(_05977_),
    .Y(_00008_)
  );
  NAND _14257_ (
    .A(\memory[10][1] ),
    .B(_05361_),
    .Y(_05978_)
  );
  OR _14258_ (
    .A(\memory[10][1] ),
    .B(_01538_),
    .Y(_05979_)
  );
  OR _14259_ (
    .A(\data_i[25] ),
    .B(_01539_),
    .Y(_05980_)
  );
  NAND _14260_ (
    .A(_05979_),
    .B(_05980_),
    .Y(_05982_)
  );
  NAND _14261_ (
    .A(_01528_),
    .B(_05982_),
    .Y(_05983_)
  );
  OR _14262_ (
    .A(\data_i[17] ),
    .B(_01528_),
    .Y(_05984_)
  );
  AND _14263_ (
    .A(_05983_),
    .B(_05984_),
    .Y(_05985_)
  );
  NAND _14264_ (
    .A(\data_i[9] ),
    .B(_01495_),
    .Y(_05986_)
  );
  AND _14265_ (
    .A(_01579_),
    .B(_05986_),
    .Y(_05987_)
  );
  NAND _14266_ (
    .A(_01496_),
    .B(_05985_),
    .Y(_05988_)
  );
  NAND _14267_ (
    .A(_05987_),
    .B(_05988_),
    .Y(_05989_)
  );
  OR _14268_ (
    .A(\data_i[1] ),
    .B(_01579_),
    .Y(_05990_)
  );
  AND _14269_ (
    .A(MemWrite_i),
    .B(_05990_),
    .Y(_05991_)
  );
  NAND _14270_ (
    .A(_05989_),
    .B(_05991_),
    .Y(_05993_)
  );
  NAND _14271_ (
    .A(_05978_),
    .B(_05993_),
    .Y(_00009_)
  );
  NAND _14272_ (
    .A(\memory[10][2] ),
    .B(_05361_),
    .Y(_05994_)
  );
  OR _14273_ (
    .A(\memory[10][2] ),
    .B(_01538_),
    .Y(_05995_)
  );
  OR _14274_ (
    .A(\data_i[26] ),
    .B(_01539_),
    .Y(_05996_)
  );
  NAND _14275_ (
    .A(_05995_),
    .B(_05996_),
    .Y(_05997_)
  );
  NAND _14276_ (
    .A(_01528_),
    .B(_05997_),
    .Y(_05998_)
  );
  OR _14277_ (
    .A(\data_i[18] ),
    .B(_01528_),
    .Y(_05999_)
  );
  AND _14278_ (
    .A(_05998_),
    .B(_05999_),
    .Y(_06000_)
  );
  NAND _14279_ (
    .A(\data_i[10] ),
    .B(_01495_),
    .Y(_06001_)
  );
  AND _14280_ (
    .A(_01579_),
    .B(_06001_),
    .Y(_06003_)
  );
  NAND _14281_ (
    .A(_01496_),
    .B(_06000_),
    .Y(_06004_)
  );
  NAND _14282_ (
    .A(_06003_),
    .B(_06004_),
    .Y(_06005_)
  );
  OR _14283_ (
    .A(\data_i[2] ),
    .B(_01579_),
    .Y(_06006_)
  );
  AND _14284_ (
    .A(MemWrite_i),
    .B(_06006_),
    .Y(_06007_)
  );
  NAND _14285_ (
    .A(_06005_),
    .B(_06007_),
    .Y(_06008_)
  );
  NAND _14286_ (
    .A(_05994_),
    .B(_06008_),
    .Y(_00010_)
  );
  NAND _14287_ (
    .A(\memory[10][3] ),
    .B(_05361_),
    .Y(_06009_)
  );
  OR _14288_ (
    .A(\memory[10][3] ),
    .B(_01538_),
    .Y(_06010_)
  );
  OR _14289_ (
    .A(\data_i[27] ),
    .B(_01539_),
    .Y(_06011_)
  );
  NAND _14290_ (
    .A(_06010_),
    .B(_06011_),
    .Y(_06013_)
  );
  NAND _14291_ (
    .A(_01528_),
    .B(_06013_),
    .Y(_06014_)
  );
  OR _14292_ (
    .A(\data_i[19] ),
    .B(_01528_),
    .Y(_06015_)
  );
  AND _14293_ (
    .A(_06014_),
    .B(_06015_),
    .Y(_06016_)
  );
  NAND _14294_ (
    .A(\data_i[11] ),
    .B(_01495_),
    .Y(_06017_)
  );
  AND _14295_ (
    .A(_01579_),
    .B(_06017_),
    .Y(_06018_)
  );
  NAND _14296_ (
    .A(_01496_),
    .B(_06016_),
    .Y(_06019_)
  );
  NAND _14297_ (
    .A(_06018_),
    .B(_06019_),
    .Y(_06020_)
  );
  OR _14298_ (
    .A(\data_i[3] ),
    .B(_01579_),
    .Y(_06021_)
  );
  AND _14299_ (
    .A(MemWrite_i),
    .B(_06021_),
    .Y(_06022_)
  );
  NAND _14300_ (
    .A(_06020_),
    .B(_06022_),
    .Y(_06024_)
  );
  NAND _14301_ (
    .A(_06009_),
    .B(_06024_),
    .Y(_00011_)
  );
  NAND _14302_ (
    .A(\memory[10][4] ),
    .B(_05361_),
    .Y(_06025_)
  );
  OR _14303_ (
    .A(\memory[10][4] ),
    .B(_01538_),
    .Y(_06026_)
  );
  OR _14304_ (
    .A(\data_i[28] ),
    .B(_01539_),
    .Y(_06027_)
  );
  NAND _14305_ (
    .A(_06026_),
    .B(_06027_),
    .Y(_06028_)
  );
  NAND _14306_ (
    .A(_01528_),
    .B(_06028_),
    .Y(_06029_)
  );
  OR _14307_ (
    .A(\data_i[20] ),
    .B(_01528_),
    .Y(_06030_)
  );
  AND _14308_ (
    .A(_06029_),
    .B(_06030_),
    .Y(_06031_)
  );
  NAND _14309_ (
    .A(\data_i[12] ),
    .B(_01495_),
    .Y(_06032_)
  );
  AND _14310_ (
    .A(_01579_),
    .B(_06032_),
    .Y(_06034_)
  );
  NAND _14311_ (
    .A(_01496_),
    .B(_06031_),
    .Y(_06035_)
  );
  NAND _14312_ (
    .A(_06034_),
    .B(_06035_),
    .Y(_06036_)
  );
  OR _14313_ (
    .A(\data_i[4] ),
    .B(_01579_),
    .Y(_06037_)
  );
  AND _14314_ (
    .A(MemWrite_i),
    .B(_06037_),
    .Y(_06038_)
  );
  NAND _14315_ (
    .A(_06036_),
    .B(_06038_),
    .Y(_06039_)
  );
  NAND _14316_ (
    .A(_06025_),
    .B(_06039_),
    .Y(_00012_)
  );
  NAND _14317_ (
    .A(\memory[10][5] ),
    .B(_05361_),
    .Y(_06040_)
  );
  OR _14318_ (
    .A(\memory[10][5] ),
    .B(_01538_),
    .Y(_06041_)
  );
  OR _14319_ (
    .A(\data_i[29] ),
    .B(_01539_),
    .Y(_06042_)
  );
  NAND _14320_ (
    .A(_06041_),
    .B(_06042_),
    .Y(_06044_)
  );
  NAND _14321_ (
    .A(_01528_),
    .B(_06044_),
    .Y(_06045_)
  );
  OR _14322_ (
    .A(\data_i[21] ),
    .B(_01528_),
    .Y(_06046_)
  );
  AND _14323_ (
    .A(_06045_),
    .B(_06046_),
    .Y(_06047_)
  );
  NAND _14324_ (
    .A(\data_i[13] ),
    .B(_01495_),
    .Y(_06048_)
  );
  AND _14325_ (
    .A(_01579_),
    .B(_06048_),
    .Y(_06049_)
  );
  NAND _14326_ (
    .A(_01496_),
    .B(_06047_),
    .Y(_06050_)
  );
  NAND _14327_ (
    .A(_06049_),
    .B(_06050_),
    .Y(_06051_)
  );
  OR _14328_ (
    .A(\data_i[5] ),
    .B(_01579_),
    .Y(_06052_)
  );
  AND _14329_ (
    .A(MemWrite_i),
    .B(_06052_),
    .Y(_06053_)
  );
  NAND _14330_ (
    .A(_06051_),
    .B(_06053_),
    .Y(_06055_)
  );
  NAND _14331_ (
    .A(_06040_),
    .B(_06055_),
    .Y(_00013_)
  );
  NAND _14332_ (
    .A(\memory[10][6] ),
    .B(_05361_),
    .Y(_06056_)
  );
  OR _14333_ (
    .A(\memory[10][6] ),
    .B(_01538_),
    .Y(_06057_)
  );
  OR _14334_ (
    .A(\data_i[30] ),
    .B(_01539_),
    .Y(_06058_)
  );
  NAND _14335_ (
    .A(_06057_),
    .B(_06058_),
    .Y(_06059_)
  );
  NAND _14336_ (
    .A(_01528_),
    .B(_06059_),
    .Y(_06060_)
  );
  OR _14337_ (
    .A(\data_i[22] ),
    .B(_01528_),
    .Y(_06061_)
  );
  AND _14338_ (
    .A(_06060_),
    .B(_06061_),
    .Y(_06062_)
  );
  NAND _14339_ (
    .A(\data_i[14] ),
    .B(_01495_),
    .Y(_06063_)
  );
  AND _14340_ (
    .A(_01579_),
    .B(_06063_),
    .Y(_06065_)
  );
  NAND _14341_ (
    .A(_01496_),
    .B(_06062_),
    .Y(_06066_)
  );
  NAND _14342_ (
    .A(_06065_),
    .B(_06066_),
    .Y(_06067_)
  );
  OR _14343_ (
    .A(\data_i[6] ),
    .B(_01579_),
    .Y(_06068_)
  );
  AND _14344_ (
    .A(MemWrite_i),
    .B(_06068_),
    .Y(_06069_)
  );
  NAND _14345_ (
    .A(_06067_),
    .B(_06069_),
    .Y(_06070_)
  );
  NAND _14346_ (
    .A(_06056_),
    .B(_06070_),
    .Y(_00014_)
  );
  NAND _14347_ (
    .A(\memory[10][7] ),
    .B(_05361_),
    .Y(_06071_)
  );
  OR _14348_ (
    .A(\memory[10][7] ),
    .B(_01538_),
    .Y(_06072_)
  );
  OR _14349_ (
    .A(\data_i[31] ),
    .B(_01539_),
    .Y(_06073_)
  );
  NAND _14350_ (
    .A(_06072_),
    .B(_06073_),
    .Y(_06075_)
  );
  NAND _14351_ (
    .A(_01528_),
    .B(_06075_),
    .Y(_06076_)
  );
  OR _14352_ (
    .A(\data_i[23] ),
    .B(_01528_),
    .Y(_06077_)
  );
  AND _14353_ (
    .A(_06076_),
    .B(_06077_),
    .Y(_06078_)
  );
  NAND _14354_ (
    .A(\data_i[15] ),
    .B(_01495_),
    .Y(_06079_)
  );
  AND _14355_ (
    .A(_01579_),
    .B(_06079_),
    .Y(_06080_)
  );
  NAND _14356_ (
    .A(_01496_),
    .B(_06078_),
    .Y(_06081_)
  );
  NAND _14357_ (
    .A(_06080_),
    .B(_06081_),
    .Y(_06082_)
  );
  OR _14358_ (
    .A(\data_i[7] ),
    .B(_01579_),
    .Y(_06083_)
  );
  AND _14359_ (
    .A(MemWrite_i),
    .B(_06083_),
    .Y(_06084_)
  );
  NAND _14360_ (
    .A(_06082_),
    .B(_06084_),
    .Y(_06086_)
  );
  NAND _14361_ (
    .A(_06071_),
    .B(_06086_),
    .Y(_00015_)
  );
  NAND _14362_ (
    .A(\memory[9][0] ),
    .B(_05361_),
    .Y(_06087_)
  );
  OR _14363_ (
    .A(\memory[9][0] ),
    .B(_01517_),
    .Y(_06088_)
  );
  OR _14364_ (
    .A(\data_i[24] ),
    .B(_01518_),
    .Y(_06089_)
  );
  NAND _14365_ (
    .A(_06088_),
    .B(_06089_),
    .Y(_06090_)
  );
  NAND _14366_ (
    .A(_01539_),
    .B(_06090_),
    .Y(_06091_)
  );
  OR _14367_ (
    .A(\data_i[16] ),
    .B(_01539_),
    .Y(_06092_)
  );
  AND _14368_ (
    .A(_06091_),
    .B(_06092_),
    .Y(_06093_)
  );
  NAND _14369_ (
    .A(\data_i[8] ),
    .B(_01527_),
    .Y(_06094_)
  );
  AND _14370_ (
    .A(_01496_),
    .B(_06094_),
    .Y(_06096_)
  );
  NAND _14371_ (
    .A(_01528_),
    .B(_06093_),
    .Y(_06097_)
  );
  NAND _14372_ (
    .A(_06096_),
    .B(_06097_),
    .Y(_06098_)
  );
  OR _14373_ (
    .A(\data_i[0] ),
    .B(_01496_),
    .Y(_06099_)
  );
  AND _14374_ (
    .A(MemWrite_i),
    .B(_06099_),
    .Y(_06100_)
  );
  NAND _14375_ (
    .A(_06098_),
    .B(_06100_),
    .Y(_06101_)
  );
  NAND _14376_ (
    .A(_06087_),
    .B(_06101_),
    .Y(_00248_)
  );
  NAND _14377_ (
    .A(\memory[9][1] ),
    .B(_05361_),
    .Y(_06102_)
  );
  OR _14378_ (
    .A(\memory[9][1] ),
    .B(_01517_),
    .Y(_06103_)
  );
  OR _14379_ (
    .A(\data_i[25] ),
    .B(_01518_),
    .Y(_06104_)
  );
  NAND _14380_ (
    .A(_06103_),
    .B(_06104_),
    .Y(_06106_)
  );
  NAND _14381_ (
    .A(_01539_),
    .B(_06106_),
    .Y(_06107_)
  );
  OR _14382_ (
    .A(\data_i[17] ),
    .B(_01539_),
    .Y(_06108_)
  );
  AND _14383_ (
    .A(_06107_),
    .B(_06108_),
    .Y(_06109_)
  );
  NAND _14384_ (
    .A(\data_i[9] ),
    .B(_01527_),
    .Y(_06110_)
  );
  AND _14385_ (
    .A(_01496_),
    .B(_06110_),
    .Y(_06111_)
  );
  NAND _14386_ (
    .A(_01528_),
    .B(_06109_),
    .Y(_06112_)
  );
  NAND _14387_ (
    .A(_06111_),
    .B(_06112_),
    .Y(_06113_)
  );
  OR _14388_ (
    .A(\data_i[1] ),
    .B(_01496_),
    .Y(_06114_)
  );
  AND _14389_ (
    .A(MemWrite_i),
    .B(_06114_),
    .Y(_06115_)
  );
  NAND _14390_ (
    .A(_06113_),
    .B(_06115_),
    .Y(_06117_)
  );
  NAND _14391_ (
    .A(_06102_),
    .B(_06117_),
    .Y(_00249_)
  );
  NAND _14392_ (
    .A(\memory[9][2] ),
    .B(_05361_),
    .Y(_06118_)
  );
  OR _14393_ (
    .A(\memory[9][2] ),
    .B(_01517_),
    .Y(_06119_)
  );
  OR _14394_ (
    .A(\data_i[26] ),
    .B(_01518_),
    .Y(_06120_)
  );
  NAND _14395_ (
    .A(_06119_),
    .B(_06120_),
    .Y(_06121_)
  );
  NAND _14396_ (
    .A(_01539_),
    .B(_06121_),
    .Y(_06122_)
  );
  OR _14397_ (
    .A(\data_i[18] ),
    .B(_01539_),
    .Y(_06123_)
  );
  AND _14398_ (
    .A(_06122_),
    .B(_06123_),
    .Y(_06124_)
  );
  NAND _14399_ (
    .A(\data_i[10] ),
    .B(_01527_),
    .Y(_06125_)
  );
  AND _14400_ (
    .A(_01496_),
    .B(_06125_),
    .Y(_06127_)
  );
  NAND _14401_ (
    .A(_01528_),
    .B(_06124_),
    .Y(_06128_)
  );
  NAND _14402_ (
    .A(_06127_),
    .B(_06128_),
    .Y(_06129_)
  );
  OR _14403_ (
    .A(\data_i[2] ),
    .B(_01496_),
    .Y(_06130_)
  );
  AND _14404_ (
    .A(MemWrite_i),
    .B(_06130_),
    .Y(_06131_)
  );
  NAND _14405_ (
    .A(_06129_),
    .B(_06131_),
    .Y(_06132_)
  );
  NAND _14406_ (
    .A(_06118_),
    .B(_06132_),
    .Y(_00250_)
  );
  NAND _14407_ (
    .A(\memory[9][3] ),
    .B(_05361_),
    .Y(_06133_)
  );
  OR _14408_ (
    .A(\memory[9][3] ),
    .B(_01517_),
    .Y(_06134_)
  );
  OR _14409_ (
    .A(\data_i[27] ),
    .B(_01518_),
    .Y(_06135_)
  );
  NAND _14410_ (
    .A(_06134_),
    .B(_06135_),
    .Y(_06137_)
  );
  NAND _14411_ (
    .A(_01539_),
    .B(_06137_),
    .Y(_06138_)
  );
  OR _14412_ (
    .A(\data_i[19] ),
    .B(_01539_),
    .Y(_06139_)
  );
  AND _14413_ (
    .A(_06138_),
    .B(_06139_),
    .Y(_06140_)
  );
  NAND _14414_ (
    .A(\data_i[11] ),
    .B(_01527_),
    .Y(_06141_)
  );
  AND _14415_ (
    .A(_01496_),
    .B(_06141_),
    .Y(_06142_)
  );
  NAND _14416_ (
    .A(_01528_),
    .B(_06140_),
    .Y(_06143_)
  );
  NAND _14417_ (
    .A(_06142_),
    .B(_06143_),
    .Y(_06144_)
  );
  OR _14418_ (
    .A(\data_i[3] ),
    .B(_01496_),
    .Y(_06145_)
  );
  AND _14419_ (
    .A(MemWrite_i),
    .B(_06145_),
    .Y(_06146_)
  );
  NAND _14420_ (
    .A(_06144_),
    .B(_06146_),
    .Y(_06148_)
  );
  NAND _14421_ (
    .A(_06133_),
    .B(_06148_),
    .Y(_00251_)
  );
  NAND _14422_ (
    .A(\memory[9][4] ),
    .B(_05361_),
    .Y(_06149_)
  );
  OR _14423_ (
    .A(\memory[9][4] ),
    .B(_01517_),
    .Y(_06150_)
  );
  OR _14424_ (
    .A(\data_i[28] ),
    .B(_01518_),
    .Y(_06151_)
  );
  NAND _14425_ (
    .A(_06150_),
    .B(_06151_),
    .Y(_06152_)
  );
  NAND _14426_ (
    .A(_01539_),
    .B(_06152_),
    .Y(_06153_)
  );
  OR _14427_ (
    .A(\data_i[20] ),
    .B(_01539_),
    .Y(_06154_)
  );
  AND _14428_ (
    .A(_06153_),
    .B(_06154_),
    .Y(_06155_)
  );
  NAND _14429_ (
    .A(\data_i[12] ),
    .B(_01527_),
    .Y(_06156_)
  );
  AND _14430_ (
    .A(_01496_),
    .B(_06156_),
    .Y(_06158_)
  );
  NAND _14431_ (
    .A(_01528_),
    .B(_06155_),
    .Y(_06159_)
  );
  NAND _14432_ (
    .A(_06158_),
    .B(_06159_),
    .Y(_06160_)
  );
  OR _14433_ (
    .A(\data_i[4] ),
    .B(_01496_),
    .Y(_06161_)
  );
  AND _14434_ (
    .A(MemWrite_i),
    .B(_06161_),
    .Y(_06162_)
  );
  NAND _14435_ (
    .A(_06160_),
    .B(_06162_),
    .Y(_06163_)
  );
  NAND _14436_ (
    .A(_06149_),
    .B(_06163_),
    .Y(_00252_)
  );
  NAND _14437_ (
    .A(\memory[9][5] ),
    .B(_05361_),
    .Y(_06164_)
  );
  OR _14438_ (
    .A(\memory[9][5] ),
    .B(_01517_),
    .Y(_06165_)
  );
  OR _14439_ (
    .A(\data_i[29] ),
    .B(_01518_),
    .Y(_06166_)
  );
  NAND _14440_ (
    .A(_06165_),
    .B(_06166_),
    .Y(_06168_)
  );
  NAND _14441_ (
    .A(_01539_),
    .B(_06168_),
    .Y(_06169_)
  );
  OR _14442_ (
    .A(\data_i[21] ),
    .B(_01539_),
    .Y(_06170_)
  );
  AND _14443_ (
    .A(_06169_),
    .B(_06170_),
    .Y(_06171_)
  );
  NAND _14444_ (
    .A(\data_i[13] ),
    .B(_01527_),
    .Y(_06172_)
  );
  AND _14445_ (
    .A(_01496_),
    .B(_06172_),
    .Y(_06173_)
  );
  NAND _14446_ (
    .A(_01528_),
    .B(_06171_),
    .Y(_06174_)
  );
  NAND _14447_ (
    .A(_06173_),
    .B(_06174_),
    .Y(_06175_)
  );
  OR _14448_ (
    .A(\data_i[5] ),
    .B(_01496_),
    .Y(_06176_)
  );
  AND _14449_ (
    .A(MemWrite_i),
    .B(_06176_),
    .Y(_06177_)
  );
  NAND _14450_ (
    .A(_06175_),
    .B(_06177_),
    .Y(_06179_)
  );
  NAND _14451_ (
    .A(_06164_),
    .B(_06179_),
    .Y(_00253_)
  );
  NAND _14452_ (
    .A(\memory[9][6] ),
    .B(_05361_),
    .Y(_06180_)
  );
  OR _14453_ (
    .A(\memory[9][6] ),
    .B(_01517_),
    .Y(_06181_)
  );
  OR _14454_ (
    .A(\data_i[30] ),
    .B(_01518_),
    .Y(_06182_)
  );
  NAND _14455_ (
    .A(_06181_),
    .B(_06182_),
    .Y(_06183_)
  );
  NAND _14456_ (
    .A(_01539_),
    .B(_06183_),
    .Y(_06184_)
  );
  OR _14457_ (
    .A(\data_i[22] ),
    .B(_01539_),
    .Y(_06185_)
  );
  AND _14458_ (
    .A(_06184_),
    .B(_06185_),
    .Y(_06186_)
  );
  NAND _14459_ (
    .A(\data_i[14] ),
    .B(_01527_),
    .Y(_06187_)
  );
  AND _14460_ (
    .A(_01496_),
    .B(_06187_),
    .Y(_06189_)
  );
  NAND _14461_ (
    .A(_01528_),
    .B(_06186_),
    .Y(_06190_)
  );
  NAND _14462_ (
    .A(_06189_),
    .B(_06190_),
    .Y(_06191_)
  );
  OR _14463_ (
    .A(\data_i[6] ),
    .B(_01496_),
    .Y(_06192_)
  );
  AND _14464_ (
    .A(MemWrite_i),
    .B(_06192_),
    .Y(_06193_)
  );
  NAND _14465_ (
    .A(_06191_),
    .B(_06193_),
    .Y(_06194_)
  );
  NAND _14466_ (
    .A(_06180_),
    .B(_06194_),
    .Y(_00254_)
  );
  NAND _14467_ (
    .A(\memory[9][7] ),
    .B(_05361_),
    .Y(_06195_)
  );
  OR _14468_ (
    .A(\memory[9][7] ),
    .B(_01517_),
    .Y(_06196_)
  );
  OR _14469_ (
    .A(\data_i[31] ),
    .B(_01518_),
    .Y(_06197_)
  );
  NAND _14470_ (
    .A(_06196_),
    .B(_06197_),
    .Y(_06199_)
  );
  NAND _14471_ (
    .A(_01539_),
    .B(_06199_),
    .Y(_06200_)
  );
  OR _14472_ (
    .A(\data_i[23] ),
    .B(_01539_),
    .Y(_06201_)
  );
  AND _14473_ (
    .A(_06200_),
    .B(_06201_),
    .Y(_06202_)
  );
  NAND _14474_ (
    .A(\data_i[15] ),
    .B(_01527_),
    .Y(_06203_)
  );
  AND _14475_ (
    .A(_01496_),
    .B(_06203_),
    .Y(_06204_)
  );
  NAND _14476_ (
    .A(_01528_),
    .B(_06202_),
    .Y(_06205_)
  );
  NAND _14477_ (
    .A(_06204_),
    .B(_06205_),
    .Y(_06206_)
  );
  OR _14478_ (
    .A(\data_i[7] ),
    .B(_01496_),
    .Y(_06207_)
  );
  AND _14479_ (
    .A(MemWrite_i),
    .B(_06207_),
    .Y(_06208_)
  );
  NAND _14480_ (
    .A(_06206_),
    .B(_06208_),
    .Y(_06210_)
  );
  NAND _14481_ (
    .A(_06195_),
    .B(_06210_),
    .Y(_00255_)
  );
  NAND _14482_ (
    .A(\memory[8][0] ),
    .B(_05361_),
    .Y(_06211_)
  );
  OR _14483_ (
    .A(\memory[8][0] ),
    .B(_01585_),
    .Y(_06212_)
  );
  OR _14484_ (
    .A(\data_i[24] ),
    .B(_01586_),
    .Y(_06213_)
  );
  NAND _14485_ (
    .A(_06212_),
    .B(_06213_),
    .Y(_06214_)
  );
  NAND _14486_ (
    .A(_01518_),
    .B(_06214_),
    .Y(_06215_)
  );
  OR _14487_ (
    .A(\data_i[16] ),
    .B(_01518_),
    .Y(_06216_)
  );
  AND _14488_ (
    .A(_06215_),
    .B(_06216_),
    .Y(_06217_)
  );
  NAND _14489_ (
    .A(\data_i[8] ),
    .B(_01538_),
    .Y(_06218_)
  );
  AND _14490_ (
    .A(_01528_),
    .B(_06218_),
    .Y(_06220_)
  );
  NAND _14491_ (
    .A(_01539_),
    .B(_06217_),
    .Y(_06221_)
  );
  NAND _14492_ (
    .A(_06220_),
    .B(_06221_),
    .Y(_06222_)
  );
  OR _14493_ (
    .A(\data_i[0] ),
    .B(_01528_),
    .Y(_06223_)
  );
  AND _14494_ (
    .A(MemWrite_i),
    .B(_06223_),
    .Y(_06224_)
  );
  NAND _14495_ (
    .A(_06222_),
    .B(_06224_),
    .Y(_06225_)
  );
  NAND _14496_ (
    .A(_06211_),
    .B(_06225_),
    .Y(_00240_)
  );
  NAND _14497_ (
    .A(\memory[8][1] ),
    .B(_05361_),
    .Y(_06226_)
  );
  OR _14498_ (
    .A(\memory[8][1] ),
    .B(_01585_),
    .Y(_06227_)
  );
  OR _14499_ (
    .A(\data_i[25] ),
    .B(_01586_),
    .Y(_06228_)
  );
  NAND _14500_ (
    .A(_06227_),
    .B(_06228_),
    .Y(_06230_)
  );
  NAND _14501_ (
    .A(_01518_),
    .B(_06230_),
    .Y(_06231_)
  );
  OR _14502_ (
    .A(\data_i[17] ),
    .B(_01518_),
    .Y(_06232_)
  );
  AND _14503_ (
    .A(_06231_),
    .B(_06232_),
    .Y(_06233_)
  );
  NAND _14504_ (
    .A(\data_i[9] ),
    .B(_01538_),
    .Y(_06234_)
  );
  AND _14505_ (
    .A(_01528_),
    .B(_06234_),
    .Y(_06235_)
  );
  NAND _14506_ (
    .A(_01539_),
    .B(_06233_),
    .Y(_06236_)
  );
  NAND _14507_ (
    .A(_06235_),
    .B(_06236_),
    .Y(_06237_)
  );
  OR _14508_ (
    .A(\data_i[1] ),
    .B(_01528_),
    .Y(_06238_)
  );
  AND _14509_ (
    .A(MemWrite_i),
    .B(_06238_),
    .Y(_06239_)
  );
  NAND _14510_ (
    .A(_06237_),
    .B(_06239_),
    .Y(_06241_)
  );
  NAND _14511_ (
    .A(_06226_),
    .B(_06241_),
    .Y(_00241_)
  );
  NAND _14512_ (
    .A(\memory[8][2] ),
    .B(_05361_),
    .Y(_06242_)
  );
  OR _14513_ (
    .A(\memory[8][2] ),
    .B(_01585_),
    .Y(_06243_)
  );
  OR _14514_ (
    .A(\data_i[26] ),
    .B(_01586_),
    .Y(_06244_)
  );
  NAND _14515_ (
    .A(_06243_),
    .B(_06244_),
    .Y(_06245_)
  );
  NAND _14516_ (
    .A(_01518_),
    .B(_06245_),
    .Y(_06246_)
  );
  OR _14517_ (
    .A(\data_i[18] ),
    .B(_01518_),
    .Y(_06247_)
  );
  AND _14518_ (
    .A(_06246_),
    .B(_06247_),
    .Y(_06248_)
  );
  NAND _14519_ (
    .A(\data_i[10] ),
    .B(_01538_),
    .Y(_06249_)
  );
  AND _14520_ (
    .A(_01528_),
    .B(_06249_),
    .Y(_06251_)
  );
  NAND _14521_ (
    .A(_01539_),
    .B(_06248_),
    .Y(_06252_)
  );
  NAND _14522_ (
    .A(_06251_),
    .B(_06252_),
    .Y(_06253_)
  );
  OR _14523_ (
    .A(\data_i[2] ),
    .B(_01528_),
    .Y(_06254_)
  );
  AND _14524_ (
    .A(MemWrite_i),
    .B(_06254_),
    .Y(_06255_)
  );
  NAND _14525_ (
    .A(_06253_),
    .B(_06255_),
    .Y(_06256_)
  );
  NAND _14526_ (
    .A(_06242_),
    .B(_06256_),
    .Y(_00242_)
  );
  NAND _14527_ (
    .A(\memory[8][3] ),
    .B(_05361_),
    .Y(_06257_)
  );
  OR _14528_ (
    .A(\memory[8][3] ),
    .B(_01585_),
    .Y(_06258_)
  );
  OR _14529_ (
    .A(\data_i[27] ),
    .B(_01586_),
    .Y(_06259_)
  );
  NAND _14530_ (
    .A(_06258_),
    .B(_06259_),
    .Y(_06261_)
  );
  NAND _14531_ (
    .A(_01518_),
    .B(_06261_),
    .Y(_06262_)
  );
  OR _14532_ (
    .A(\data_i[19] ),
    .B(_01518_),
    .Y(_06263_)
  );
  AND _14533_ (
    .A(_06262_),
    .B(_06263_),
    .Y(_06264_)
  );
  NAND _14534_ (
    .A(\data_i[11] ),
    .B(_01538_),
    .Y(_06265_)
  );
  AND _14535_ (
    .A(_01528_),
    .B(_06265_),
    .Y(_06266_)
  );
  NAND _14536_ (
    .A(_01539_),
    .B(_06264_),
    .Y(_06267_)
  );
  NAND _14537_ (
    .A(_06266_),
    .B(_06267_),
    .Y(_06268_)
  );
  OR _14538_ (
    .A(\data_i[3] ),
    .B(_01528_),
    .Y(_06269_)
  );
  AND _14539_ (
    .A(MemWrite_i),
    .B(_06269_),
    .Y(_06270_)
  );
  NAND _14540_ (
    .A(_06268_),
    .B(_06270_),
    .Y(_06272_)
  );
  NAND _14541_ (
    .A(_06257_),
    .B(_06272_),
    .Y(_00243_)
  );
  NAND _14542_ (
    .A(\memory[8][4] ),
    .B(_05361_),
    .Y(_06273_)
  );
  OR _14543_ (
    .A(\memory[8][4] ),
    .B(_01585_),
    .Y(_06274_)
  );
  OR _14544_ (
    .A(\data_i[28] ),
    .B(_01586_),
    .Y(_06275_)
  );
  NAND _14545_ (
    .A(_06274_),
    .B(_06275_),
    .Y(_06276_)
  );
  NAND _14546_ (
    .A(_01518_),
    .B(_06276_),
    .Y(_06277_)
  );
  OR _14547_ (
    .A(\data_i[20] ),
    .B(_01518_),
    .Y(_06278_)
  );
  AND _14548_ (
    .A(_06277_),
    .B(_06278_),
    .Y(_06279_)
  );
  NAND _14549_ (
    .A(\data_i[12] ),
    .B(_01538_),
    .Y(_06280_)
  );
  AND _14550_ (
    .A(_01528_),
    .B(_06280_),
    .Y(_06282_)
  );
  NAND _14551_ (
    .A(_01539_),
    .B(_06279_),
    .Y(_06283_)
  );
  NAND _14552_ (
    .A(_06282_),
    .B(_06283_),
    .Y(_06284_)
  );
  OR _14553_ (
    .A(\data_i[4] ),
    .B(_01528_),
    .Y(_06285_)
  );
  AND _14554_ (
    .A(MemWrite_i),
    .B(_06285_),
    .Y(_06286_)
  );
  NAND _14555_ (
    .A(_06284_),
    .B(_06286_),
    .Y(_06287_)
  );
  NAND _14556_ (
    .A(_06273_),
    .B(_06287_),
    .Y(_00244_)
  );
  NAND _14557_ (
    .A(\memory[8][5] ),
    .B(_05361_),
    .Y(_06288_)
  );
  OR _14558_ (
    .A(\memory[8][5] ),
    .B(_01585_),
    .Y(_06289_)
  );
  OR _14559_ (
    .A(\data_i[29] ),
    .B(_01586_),
    .Y(_06290_)
  );
  NAND _14560_ (
    .A(_06289_),
    .B(_06290_),
    .Y(_06292_)
  );
  NAND _14561_ (
    .A(_01518_),
    .B(_06292_),
    .Y(_06293_)
  );
  OR _14562_ (
    .A(\data_i[21] ),
    .B(_01518_),
    .Y(_06294_)
  );
  AND _14563_ (
    .A(_06293_),
    .B(_06294_),
    .Y(_06295_)
  );
  NAND _14564_ (
    .A(\data_i[13] ),
    .B(_01538_),
    .Y(_06296_)
  );
  AND _14565_ (
    .A(_01528_),
    .B(_06296_),
    .Y(_06297_)
  );
  NAND _14566_ (
    .A(_01539_),
    .B(_06295_),
    .Y(_06298_)
  );
  NAND _14567_ (
    .A(_06297_),
    .B(_06298_),
    .Y(_06299_)
  );
  OR _14568_ (
    .A(\data_i[5] ),
    .B(_01528_),
    .Y(_06300_)
  );
  AND _14569_ (
    .A(MemWrite_i),
    .B(_06300_),
    .Y(_06301_)
  );
  NAND _14570_ (
    .A(_06299_),
    .B(_06301_),
    .Y(_06303_)
  );
  NAND _14571_ (
    .A(_06288_),
    .B(_06303_),
    .Y(_00245_)
  );
  NAND _14572_ (
    .A(\memory[8][6] ),
    .B(_05361_),
    .Y(_06304_)
  );
  OR _14573_ (
    .A(\memory[8][6] ),
    .B(_01585_),
    .Y(_06305_)
  );
  OR _14574_ (
    .A(\data_i[30] ),
    .B(_01586_),
    .Y(_06306_)
  );
  NAND _14575_ (
    .A(_06305_),
    .B(_06306_),
    .Y(_06307_)
  );
  NAND _14576_ (
    .A(_01518_),
    .B(_06307_),
    .Y(_06308_)
  );
  OR _14577_ (
    .A(\data_i[22] ),
    .B(_01518_),
    .Y(_06309_)
  );
  AND _14578_ (
    .A(_06308_),
    .B(_06309_),
    .Y(_06310_)
  );
  NAND _14579_ (
    .A(\data_i[14] ),
    .B(_01538_),
    .Y(_06311_)
  );
  AND _14580_ (
    .A(_01528_),
    .B(_06311_),
    .Y(_06313_)
  );
  NAND _14581_ (
    .A(_01539_),
    .B(_06310_),
    .Y(_06314_)
  );
  NAND _14582_ (
    .A(_06313_),
    .B(_06314_),
    .Y(_06315_)
  );
  OR _14583_ (
    .A(\data_i[6] ),
    .B(_01528_),
    .Y(_06316_)
  );
  AND _14584_ (
    .A(MemWrite_i),
    .B(_06316_),
    .Y(_06317_)
  );
  NAND _14585_ (
    .A(_06315_),
    .B(_06317_),
    .Y(_06318_)
  );
  NAND _14586_ (
    .A(_06304_),
    .B(_06318_),
    .Y(_00246_)
  );
  NAND _14587_ (
    .A(\memory[8][7] ),
    .B(_05361_),
    .Y(_06319_)
  );
  OR _14588_ (
    .A(\memory[8][7] ),
    .B(_01585_),
    .Y(_06320_)
  );
  OR _14589_ (
    .A(\data_i[31] ),
    .B(_01586_),
    .Y(_06321_)
  );
  NAND _14590_ (
    .A(_06320_),
    .B(_06321_),
    .Y(_06323_)
  );
  NAND _14591_ (
    .A(_01518_),
    .B(_06323_),
    .Y(_06324_)
  );
  OR _14592_ (
    .A(\data_i[23] ),
    .B(_01518_),
    .Y(_06325_)
  );
  AND _14593_ (
    .A(_06324_),
    .B(_06325_),
    .Y(_06326_)
  );
  NAND _14594_ (
    .A(\data_i[15] ),
    .B(_01538_),
    .Y(_06327_)
  );
  AND _14595_ (
    .A(_01528_),
    .B(_06327_),
    .Y(_06328_)
  );
  NAND _14596_ (
    .A(_01539_),
    .B(_06326_),
    .Y(_06329_)
  );
  NAND _14597_ (
    .A(_06328_),
    .B(_06329_),
    .Y(_06330_)
  );
  OR _14598_ (
    .A(\data_i[7] ),
    .B(_01528_),
    .Y(_06331_)
  );
  AND _14599_ (
    .A(MemWrite_i),
    .B(_06331_),
    .Y(_06332_)
  );
  NAND _14600_ (
    .A(_06330_),
    .B(_06332_),
    .Y(_06334_)
  );
  NAND _14601_ (
    .A(_06319_),
    .B(_06334_),
    .Y(_00247_)
  );
  NAND _14602_ (
    .A(\memory[7][0] ),
    .B(_05361_),
    .Y(_06335_)
  );
  OR _14603_ (
    .A(\memory[7][0] ),
    .B(_01530_),
    .Y(_06336_)
  );
  OR _14604_ (
    .A(\data_i[24] ),
    .B(_01531_),
    .Y(_06337_)
  );
  NAND _14605_ (
    .A(_06336_),
    .B(_06337_),
    .Y(_06338_)
  );
  NAND _14606_ (
    .A(_01586_),
    .B(_06338_),
    .Y(_06339_)
  );
  OR _14607_ (
    .A(\data_i[16] ),
    .B(_01586_),
    .Y(_06340_)
  );
  AND _14608_ (
    .A(_06339_),
    .B(_06340_),
    .Y(_06341_)
  );
  NAND _14609_ (
    .A(\data_i[8] ),
    .B(_01517_),
    .Y(_06342_)
  );
  AND _14610_ (
    .A(_01539_),
    .B(_06342_),
    .Y(_06344_)
  );
  NAND _14611_ (
    .A(_01518_),
    .B(_06341_),
    .Y(_06345_)
  );
  NAND _14612_ (
    .A(_06344_),
    .B(_06345_),
    .Y(_06346_)
  );
  OR _14613_ (
    .A(\data_i[0] ),
    .B(_01539_),
    .Y(_06347_)
  );
  AND _14614_ (
    .A(MemWrite_i),
    .B(_06347_),
    .Y(_06348_)
  );
  NAND _14615_ (
    .A(_06346_),
    .B(_06348_),
    .Y(_06349_)
  );
  NAND _14616_ (
    .A(_06335_),
    .B(_06349_),
    .Y(_00232_)
  );
  NAND _14617_ (
    .A(\memory[7][1] ),
    .B(_05361_),
    .Y(_06350_)
  );
  OR _14618_ (
    .A(\memory[7][1] ),
    .B(_01530_),
    .Y(_06351_)
  );
  OR _14619_ (
    .A(\data_i[25] ),
    .B(_01531_),
    .Y(_06352_)
  );
  NAND _14620_ (
    .A(_06351_),
    .B(_06352_),
    .Y(_06354_)
  );
  NAND _14621_ (
    .A(_01586_),
    .B(_06354_),
    .Y(_06355_)
  );
  OR _14622_ (
    .A(\data_i[17] ),
    .B(_01586_),
    .Y(_06356_)
  );
  AND _14623_ (
    .A(_06355_),
    .B(_06356_),
    .Y(_06357_)
  );
  NAND _14624_ (
    .A(_01518_),
    .B(_06357_),
    .Y(_06358_)
  );
  NAND _14625_ (
    .A(\data_i[9] ),
    .B(_01517_),
    .Y(_06359_)
  );
  AND _14626_ (
    .A(_01539_),
    .B(_06359_),
    .Y(_06360_)
  );
  NAND _14627_ (
    .A(_06358_),
    .B(_06360_),
    .Y(_06361_)
  );
  OR _14628_ (
    .A(\data_i[1] ),
    .B(_01539_),
    .Y(_06362_)
  );
  AND _14629_ (
    .A(MemWrite_i),
    .B(_06362_),
    .Y(_06363_)
  );
  NAND _14630_ (
    .A(_06361_),
    .B(_06363_),
    .Y(_06365_)
  );
  NAND _14631_ (
    .A(_06350_),
    .B(_06365_),
    .Y(_00233_)
  );
  NAND _14632_ (
    .A(\memory[7][2] ),
    .B(_05361_),
    .Y(_06366_)
  );
  OR _14633_ (
    .A(\memory[7][2] ),
    .B(_01530_),
    .Y(_06367_)
  );
  OR _14634_ (
    .A(\data_i[26] ),
    .B(_01531_),
    .Y(_06368_)
  );
  NAND _14635_ (
    .A(_06367_),
    .B(_06368_),
    .Y(_06369_)
  );
  NAND _14636_ (
    .A(_01586_),
    .B(_06369_),
    .Y(_06370_)
  );
  OR _14637_ (
    .A(\data_i[18] ),
    .B(_01586_),
    .Y(_06371_)
  );
  AND _14638_ (
    .A(_06370_),
    .B(_06371_),
    .Y(_06372_)
  );
  NAND _14639_ (
    .A(\data_i[10] ),
    .B(_01517_),
    .Y(_06373_)
  );
  AND _14640_ (
    .A(_01539_),
    .B(_06373_),
    .Y(_06375_)
  );
  NAND _14641_ (
    .A(_01518_),
    .B(_06372_),
    .Y(_06376_)
  );
  NAND _14642_ (
    .A(_06375_),
    .B(_06376_),
    .Y(_06377_)
  );
  OR _14643_ (
    .A(\data_i[2] ),
    .B(_01539_),
    .Y(_06378_)
  );
  AND _14644_ (
    .A(MemWrite_i),
    .B(_06378_),
    .Y(_06379_)
  );
  NAND _14645_ (
    .A(_06377_),
    .B(_06379_),
    .Y(_06380_)
  );
  NAND _14646_ (
    .A(_06366_),
    .B(_06380_),
    .Y(_00234_)
  );
  NAND _14647_ (
    .A(\memory[7][3] ),
    .B(_05361_),
    .Y(_06381_)
  );
  OR _14648_ (
    .A(\memory[7][3] ),
    .B(_01530_),
    .Y(_06382_)
  );
  OR _14649_ (
    .A(\data_i[27] ),
    .B(_01531_),
    .Y(_06383_)
  );
  NAND _14650_ (
    .A(_06382_),
    .B(_06383_),
    .Y(_06385_)
  );
  NAND _14651_ (
    .A(_01586_),
    .B(_06385_),
    .Y(_06386_)
  );
  OR _14652_ (
    .A(\data_i[19] ),
    .B(_01586_),
    .Y(_06387_)
  );
  AND _14653_ (
    .A(_06386_),
    .B(_06387_),
    .Y(_06388_)
  );
  NAND _14654_ (
    .A(\data_i[11] ),
    .B(_01517_),
    .Y(_06389_)
  );
  AND _14655_ (
    .A(_01539_),
    .B(_06389_),
    .Y(_06390_)
  );
  NAND _14656_ (
    .A(_01518_),
    .B(_06388_),
    .Y(_06391_)
  );
  NAND _14657_ (
    .A(_06390_),
    .B(_06391_),
    .Y(_06392_)
  );
  OR _14658_ (
    .A(\data_i[3] ),
    .B(_01539_),
    .Y(_06393_)
  );
  AND _14659_ (
    .A(MemWrite_i),
    .B(_06393_),
    .Y(_06394_)
  );
  NAND _14660_ (
    .A(_06392_),
    .B(_06394_),
    .Y(_06396_)
  );
  NAND _14661_ (
    .A(_06381_),
    .B(_06396_),
    .Y(_00235_)
  );
  NAND _14662_ (
    .A(\memory[7][4] ),
    .B(_05361_),
    .Y(_06397_)
  );
  OR _14663_ (
    .A(\memory[7][4] ),
    .B(_01530_),
    .Y(_06398_)
  );
  OR _14664_ (
    .A(\data_i[28] ),
    .B(_01531_),
    .Y(_06399_)
  );
  NAND _14665_ (
    .A(_06398_),
    .B(_06399_),
    .Y(_06400_)
  );
  NAND _14666_ (
    .A(_01586_),
    .B(_06400_),
    .Y(_06401_)
  );
  OR _14667_ (
    .A(\data_i[20] ),
    .B(_01586_),
    .Y(_06402_)
  );
  AND _14668_ (
    .A(_06401_),
    .B(_06402_),
    .Y(_06403_)
  );
  NAND _14669_ (
    .A(\data_i[12] ),
    .B(_01517_),
    .Y(_06404_)
  );
  AND _14670_ (
    .A(_01539_),
    .B(_06404_),
    .Y(_06406_)
  );
  NAND _14671_ (
    .A(_01518_),
    .B(_06403_),
    .Y(_06407_)
  );
  NAND _14672_ (
    .A(_06406_),
    .B(_06407_),
    .Y(_06408_)
  );
  OR _14673_ (
    .A(\data_i[4] ),
    .B(_01539_),
    .Y(_06409_)
  );
  AND _14674_ (
    .A(MemWrite_i),
    .B(_06409_),
    .Y(_06410_)
  );
  NAND _14675_ (
    .A(_06408_),
    .B(_06410_),
    .Y(_06411_)
  );
  NAND _14676_ (
    .A(_06397_),
    .B(_06411_),
    .Y(_00236_)
  );
  NAND _14677_ (
    .A(\memory[7][5] ),
    .B(_05361_),
    .Y(_06412_)
  );
  OR _14678_ (
    .A(\memory[7][5] ),
    .B(_01530_),
    .Y(_06413_)
  );
  OR _14679_ (
    .A(\data_i[29] ),
    .B(_01531_),
    .Y(_06414_)
  );
  NAND _14680_ (
    .A(_06413_),
    .B(_06414_),
    .Y(_06416_)
  );
  NAND _14681_ (
    .A(_01586_),
    .B(_06416_),
    .Y(_06417_)
  );
  OR _14682_ (
    .A(\data_i[21] ),
    .B(_01586_),
    .Y(_06418_)
  );
  AND _14683_ (
    .A(_06417_),
    .B(_06418_),
    .Y(_06419_)
  );
  NAND _14684_ (
    .A(\data_i[13] ),
    .B(_01517_),
    .Y(_06420_)
  );
  AND _14685_ (
    .A(_01539_),
    .B(_06420_),
    .Y(_06421_)
  );
  NAND _14686_ (
    .A(_01518_),
    .B(_06419_),
    .Y(_06422_)
  );
  NAND _14687_ (
    .A(_06421_),
    .B(_06422_),
    .Y(_06423_)
  );
  OR _14688_ (
    .A(\data_i[5] ),
    .B(_01539_),
    .Y(_06424_)
  );
  AND _14689_ (
    .A(MemWrite_i),
    .B(_06424_),
    .Y(_06425_)
  );
  NAND _14690_ (
    .A(_06423_),
    .B(_06425_),
    .Y(_06427_)
  );
  NAND _14691_ (
    .A(_06412_),
    .B(_06427_),
    .Y(_00237_)
  );
  NAND _14692_ (
    .A(\memory[7][6] ),
    .B(_05361_),
    .Y(_06428_)
  );
  OR _14693_ (
    .A(\memory[7][6] ),
    .B(_01530_),
    .Y(_06429_)
  );
  OR _14694_ (
    .A(\data_i[30] ),
    .B(_01531_),
    .Y(_06430_)
  );
  NAND _14695_ (
    .A(_06429_),
    .B(_06430_),
    .Y(_06431_)
  );
  NAND _14696_ (
    .A(_01586_),
    .B(_06431_),
    .Y(_06432_)
  );
  OR _14697_ (
    .A(\data_i[22] ),
    .B(_01586_),
    .Y(_06433_)
  );
  AND _14698_ (
    .A(_06432_),
    .B(_06433_),
    .Y(_06434_)
  );
  NAND _14699_ (
    .A(\data_i[14] ),
    .B(_01517_),
    .Y(_06435_)
  );
  AND _14700_ (
    .A(_01539_),
    .B(_06435_),
    .Y(_06437_)
  );
  NAND _14701_ (
    .A(_01518_),
    .B(_06434_),
    .Y(_06438_)
  );
  NAND _14702_ (
    .A(_06437_),
    .B(_06438_),
    .Y(_06439_)
  );
  OR _14703_ (
    .A(\data_i[6] ),
    .B(_01539_),
    .Y(_06440_)
  );
  AND _14704_ (
    .A(MemWrite_i),
    .B(_06440_),
    .Y(_06441_)
  );
  NAND _14705_ (
    .A(_06439_),
    .B(_06441_),
    .Y(_06442_)
  );
  NAND _14706_ (
    .A(_06428_),
    .B(_06442_),
    .Y(_00238_)
  );
  NAND _14707_ (
    .A(\memory[7][7] ),
    .B(_05361_),
    .Y(_06443_)
  );
  OR _14708_ (
    .A(\memory[7][7] ),
    .B(_01530_),
    .Y(_06444_)
  );
  OR _14709_ (
    .A(\data_i[31] ),
    .B(_01531_),
    .Y(_06445_)
  );
  NAND _14710_ (
    .A(_06444_),
    .B(_06445_),
    .Y(_06447_)
  );
  NAND _14711_ (
    .A(_01586_),
    .B(_06447_),
    .Y(_06448_)
  );
  OR _14712_ (
    .A(\data_i[23] ),
    .B(_01586_),
    .Y(_06449_)
  );
  AND _14713_ (
    .A(_06448_),
    .B(_06449_),
    .Y(_06450_)
  );
  NAND _14714_ (
    .A(\data_i[15] ),
    .B(_01517_),
    .Y(_06451_)
  );
  AND _14715_ (
    .A(_01539_),
    .B(_06451_),
    .Y(_06452_)
  );
  NAND _14716_ (
    .A(_01518_),
    .B(_06450_),
    .Y(_06453_)
  );
  NAND _14717_ (
    .A(_06452_),
    .B(_06453_),
    .Y(_06454_)
  );
  OR _14718_ (
    .A(\data_i[7] ),
    .B(_01539_),
    .Y(_06455_)
  );
  AND _14719_ (
    .A(MemWrite_i),
    .B(_06455_),
    .Y(_06456_)
  );
  NAND _14720_ (
    .A(_06454_),
    .B(_06456_),
    .Y(_06458_)
  );
  NAND _14721_ (
    .A(_06443_),
    .B(_06458_),
    .Y(_00239_)
  );
  NAND _14722_ (
    .A(\memory[6][0] ),
    .B(_05361_),
    .Y(_06459_)
  );
  OR _14723_ (
    .A(\memory[6][0] ),
    .B(_01513_),
    .Y(_06460_)
  );
  OR _14724_ (
    .A(\data_i[24] ),
    .B(_01514_),
    .Y(_06461_)
  );
  NAND _14725_ (
    .A(_06460_),
    .B(_06461_),
    .Y(_06462_)
  );
  NAND _14726_ (
    .A(_01531_),
    .B(_06462_),
    .Y(_06463_)
  );
  OR _14727_ (
    .A(\data_i[16] ),
    .B(_01531_),
    .Y(_06464_)
  );
  AND _14728_ (
    .A(_06463_),
    .B(_06464_),
    .Y(_06465_)
  );
  NAND _14729_ (
    .A(\data_i[8] ),
    .B(_01585_),
    .Y(_06466_)
  );
  AND _14730_ (
    .A(_01518_),
    .B(_06466_),
    .Y(_06468_)
  );
  NAND _14731_ (
    .A(_01586_),
    .B(_06465_),
    .Y(_06469_)
  );
  NAND _14732_ (
    .A(_06468_),
    .B(_06469_),
    .Y(_06470_)
  );
  OR _14733_ (
    .A(\data_i[0] ),
    .B(_01518_),
    .Y(_06471_)
  );
  AND _14734_ (
    .A(MemWrite_i),
    .B(_06471_),
    .Y(_06472_)
  );
  NAND _14735_ (
    .A(_06470_),
    .B(_06472_),
    .Y(_06473_)
  );
  NAND _14736_ (
    .A(_06459_),
    .B(_06473_),
    .Y(_00224_)
  );
  NAND _14737_ (
    .A(\memory[6][1] ),
    .B(_05361_),
    .Y(_06474_)
  );
  OR _14738_ (
    .A(\memory[6][1] ),
    .B(_01513_),
    .Y(_06475_)
  );
  OR _14739_ (
    .A(\data_i[25] ),
    .B(_01514_),
    .Y(_06476_)
  );
  NAND _14740_ (
    .A(_06475_),
    .B(_06476_),
    .Y(_06478_)
  );
  NAND _14741_ (
    .A(_01531_),
    .B(_06478_),
    .Y(_06479_)
  );
  OR _14742_ (
    .A(\data_i[17] ),
    .B(_01531_),
    .Y(_06480_)
  );
  AND _14743_ (
    .A(_06479_),
    .B(_06480_),
    .Y(_06481_)
  );
  NAND _14744_ (
    .A(\data_i[9] ),
    .B(_01585_),
    .Y(_06482_)
  );
  AND _14745_ (
    .A(_01518_),
    .B(_06482_),
    .Y(_06483_)
  );
  NAND _14746_ (
    .A(_01586_),
    .B(_06481_),
    .Y(_06484_)
  );
  NAND _14747_ (
    .A(_06483_),
    .B(_06484_),
    .Y(_06485_)
  );
  OR _14748_ (
    .A(\data_i[1] ),
    .B(_01518_),
    .Y(_06486_)
  );
  AND _14749_ (
    .A(MemWrite_i),
    .B(_06486_),
    .Y(_06487_)
  );
  NAND _14750_ (
    .A(_06485_),
    .B(_06487_),
    .Y(_06489_)
  );
  NAND _14751_ (
    .A(_06474_),
    .B(_06489_),
    .Y(_00225_)
  );
  NAND _14752_ (
    .A(\memory[6][2] ),
    .B(_05361_),
    .Y(_06490_)
  );
  OR _14753_ (
    .A(\memory[6][2] ),
    .B(_01513_),
    .Y(_06491_)
  );
  OR _14754_ (
    .A(\data_i[26] ),
    .B(_01514_),
    .Y(_06492_)
  );
  NAND _14755_ (
    .A(_06491_),
    .B(_06492_),
    .Y(_06493_)
  );
  NAND _14756_ (
    .A(_01531_),
    .B(_06493_),
    .Y(_06494_)
  );
  OR _14757_ (
    .A(\data_i[18] ),
    .B(_01531_),
    .Y(_06495_)
  );
  AND _14758_ (
    .A(_06494_),
    .B(_06495_),
    .Y(_06496_)
  );
  NAND _14759_ (
    .A(\data_i[10] ),
    .B(_01585_),
    .Y(_06497_)
  );
  AND _14760_ (
    .A(_01518_),
    .B(_06497_),
    .Y(_06499_)
  );
  NAND _14761_ (
    .A(_01586_),
    .B(_06496_),
    .Y(_06500_)
  );
  NAND _14762_ (
    .A(_06499_),
    .B(_06500_),
    .Y(_06501_)
  );
  OR _14763_ (
    .A(\data_i[2] ),
    .B(_01518_),
    .Y(_06502_)
  );
  AND _14764_ (
    .A(MemWrite_i),
    .B(_06502_),
    .Y(_06503_)
  );
  NAND _14765_ (
    .A(_06501_),
    .B(_06503_),
    .Y(_06504_)
  );
  NAND _14766_ (
    .A(_06490_),
    .B(_06504_),
    .Y(_00226_)
  );
  NAND _14767_ (
    .A(\memory[6][3] ),
    .B(_05361_),
    .Y(_06505_)
  );
  OR _14768_ (
    .A(\memory[6][3] ),
    .B(_01513_),
    .Y(_06506_)
  );
  OR _14769_ (
    .A(\data_i[27] ),
    .B(_01514_),
    .Y(_06507_)
  );
  NAND _14770_ (
    .A(_06506_),
    .B(_06507_),
    .Y(_06509_)
  );
  NAND _14771_ (
    .A(_01531_),
    .B(_06509_),
    .Y(_06510_)
  );
  OR _14772_ (
    .A(\data_i[19] ),
    .B(_01531_),
    .Y(_06511_)
  );
  AND _14773_ (
    .A(_06510_),
    .B(_06511_),
    .Y(_06512_)
  );
  NAND _14774_ (
    .A(\data_i[11] ),
    .B(_01585_),
    .Y(_06513_)
  );
  AND _14775_ (
    .A(_01518_),
    .B(_06513_),
    .Y(_06514_)
  );
  NAND _14776_ (
    .A(_01586_),
    .B(_06512_),
    .Y(_06515_)
  );
  NAND _14777_ (
    .A(_06514_),
    .B(_06515_),
    .Y(_06516_)
  );
  OR _14778_ (
    .A(\data_i[3] ),
    .B(_01518_),
    .Y(_06517_)
  );
  AND _14779_ (
    .A(MemWrite_i),
    .B(_06517_),
    .Y(_06518_)
  );
  NAND _14780_ (
    .A(_06516_),
    .B(_06518_),
    .Y(_06520_)
  );
  NAND _14781_ (
    .A(_06505_),
    .B(_06520_),
    .Y(_00227_)
  );
  NAND _14782_ (
    .A(\memory[6][4] ),
    .B(_05361_),
    .Y(_06521_)
  );
  OR _14783_ (
    .A(\memory[6][4] ),
    .B(_01513_),
    .Y(_06522_)
  );
  OR _14784_ (
    .A(\data_i[28] ),
    .B(_01514_),
    .Y(_06523_)
  );
  NAND _14785_ (
    .A(_06522_),
    .B(_06523_),
    .Y(_06524_)
  );
  NAND _14786_ (
    .A(_01531_),
    .B(_06524_),
    .Y(_06525_)
  );
  OR _14787_ (
    .A(\data_i[20] ),
    .B(_01531_),
    .Y(_06526_)
  );
  AND _14788_ (
    .A(_06525_),
    .B(_06526_),
    .Y(_06527_)
  );
  NAND _14789_ (
    .A(\data_i[12] ),
    .B(_01585_),
    .Y(_06528_)
  );
  AND _14790_ (
    .A(_01518_),
    .B(_06528_),
    .Y(_06530_)
  );
  NAND _14791_ (
    .A(_01586_),
    .B(_06527_),
    .Y(_06531_)
  );
  NAND _14792_ (
    .A(_06530_),
    .B(_06531_),
    .Y(_06532_)
  );
  OR _14793_ (
    .A(\data_i[4] ),
    .B(_01518_),
    .Y(_06533_)
  );
  AND _14794_ (
    .A(MemWrite_i),
    .B(_06533_),
    .Y(_06534_)
  );
  NAND _14795_ (
    .A(_06532_),
    .B(_06534_),
    .Y(_06535_)
  );
  NAND _14796_ (
    .A(_06521_),
    .B(_06535_),
    .Y(_00228_)
  );
  NAND _14797_ (
    .A(\memory[6][5] ),
    .B(_05361_),
    .Y(_06536_)
  );
  OR _14798_ (
    .A(\memory[6][5] ),
    .B(_01513_),
    .Y(_06537_)
  );
  OR _14799_ (
    .A(\data_i[29] ),
    .B(_01514_),
    .Y(_06538_)
  );
  NAND _14800_ (
    .A(_06537_),
    .B(_06538_),
    .Y(_06540_)
  );
  NAND _14801_ (
    .A(_01531_),
    .B(_06540_),
    .Y(_06541_)
  );
  OR _14802_ (
    .A(\data_i[21] ),
    .B(_01531_),
    .Y(_06542_)
  );
  AND _14803_ (
    .A(_06541_),
    .B(_06542_),
    .Y(_06543_)
  );
  NAND _14804_ (
    .A(\data_i[13] ),
    .B(_01585_),
    .Y(_06544_)
  );
  AND _14805_ (
    .A(_01518_),
    .B(_06544_),
    .Y(_06545_)
  );
  NAND _14806_ (
    .A(_01586_),
    .B(_06543_),
    .Y(_06546_)
  );
  NAND _14807_ (
    .A(_06545_),
    .B(_06546_),
    .Y(_06547_)
  );
  OR _14808_ (
    .A(\data_i[5] ),
    .B(_01518_),
    .Y(_06548_)
  );
  AND _14809_ (
    .A(MemWrite_i),
    .B(_06548_),
    .Y(_06549_)
  );
  NAND _14810_ (
    .A(_06547_),
    .B(_06549_),
    .Y(_06551_)
  );
  NAND _14811_ (
    .A(_06536_),
    .B(_06551_),
    .Y(_00229_)
  );
  NAND _14812_ (
    .A(\memory[6][6] ),
    .B(_05361_),
    .Y(_06552_)
  );
  OR _14813_ (
    .A(\memory[6][6] ),
    .B(_01513_),
    .Y(_06553_)
  );
  OR _14814_ (
    .A(\data_i[30] ),
    .B(_01514_),
    .Y(_06554_)
  );
  NAND _14815_ (
    .A(_06553_),
    .B(_06554_),
    .Y(_06555_)
  );
  NAND _14816_ (
    .A(_01531_),
    .B(_06555_),
    .Y(_06556_)
  );
  OR _14817_ (
    .A(\data_i[22] ),
    .B(_01531_),
    .Y(_06557_)
  );
  AND _14818_ (
    .A(_06556_),
    .B(_06557_),
    .Y(_06558_)
  );
  NAND _14819_ (
    .A(\data_i[14] ),
    .B(_01585_),
    .Y(_06559_)
  );
  AND _14820_ (
    .A(_01518_),
    .B(_06559_),
    .Y(_06561_)
  );
  NAND _14821_ (
    .A(_01586_),
    .B(_06558_),
    .Y(_06562_)
  );
  NAND _14822_ (
    .A(_06561_),
    .B(_06562_),
    .Y(_06563_)
  );
  OR _14823_ (
    .A(\data_i[6] ),
    .B(_01518_),
    .Y(_06564_)
  );
  AND _14824_ (
    .A(MemWrite_i),
    .B(_06564_),
    .Y(_06565_)
  );
  NAND _14825_ (
    .A(_06563_),
    .B(_06565_),
    .Y(_06566_)
  );
  NAND _14826_ (
    .A(_06552_),
    .B(_06566_),
    .Y(_00230_)
  );
  NAND _14827_ (
    .A(\memory[6][7] ),
    .B(_05361_),
    .Y(_06567_)
  );
  OR _14828_ (
    .A(\memory[6][7] ),
    .B(_01513_),
    .Y(_06568_)
  );
  OR _14829_ (
    .A(\data_i[31] ),
    .B(_01514_),
    .Y(_06569_)
  );
  NAND _14830_ (
    .A(_06568_),
    .B(_06569_),
    .Y(_06571_)
  );
  NAND _14831_ (
    .A(_01531_),
    .B(_06571_),
    .Y(_06572_)
  );
  OR _14832_ (
    .A(\data_i[23] ),
    .B(_01531_),
    .Y(_06573_)
  );
  AND _14833_ (
    .A(_06572_),
    .B(_06573_),
    .Y(_06574_)
  );
  NAND _14834_ (
    .A(\data_i[15] ),
    .B(_01585_),
    .Y(_06575_)
  );
  AND _14835_ (
    .A(_01518_),
    .B(_06575_),
    .Y(_06576_)
  );
  NAND _14836_ (
    .A(_01586_),
    .B(_06574_),
    .Y(_06577_)
  );
  NAND _14837_ (
    .A(_06576_),
    .B(_06577_),
    .Y(_06578_)
  );
  OR _14838_ (
    .A(\data_i[7] ),
    .B(_01518_),
    .Y(_06579_)
  );
  AND _14839_ (
    .A(MemWrite_i),
    .B(_06579_),
    .Y(_06580_)
  );
  NAND _14840_ (
    .A(_06578_),
    .B(_06580_),
    .Y(_06582_)
  );
  NAND _14841_ (
    .A(_06567_),
    .B(_06582_),
    .Y(_00231_)
  );
  NAND _14842_ (
    .A(\memory[5][0] ),
    .B(_05361_),
    .Y(_06583_)
  );
  OR _14843_ (
    .A(\memory[5][0] ),
    .B(_01453_),
    .Y(_06584_)
  );
  OR _14844_ (
    .A(\data_i[24] ),
    .B(_01454_),
    .Y(_06585_)
  );
  NAND _14845_ (
    .A(_06584_),
    .B(_06585_),
    .Y(_06586_)
  );
  NAND _14846_ (
    .A(_01514_),
    .B(_06586_),
    .Y(_06587_)
  );
  OR _14847_ (
    .A(\data_i[16] ),
    .B(_01514_),
    .Y(_06588_)
  );
  AND _14848_ (
    .A(_06587_),
    .B(_06588_),
    .Y(_06589_)
  );
  NAND _14849_ (
    .A(\data_i[8] ),
    .B(_01530_),
    .Y(_06590_)
  );
  AND _14850_ (
    .A(_01586_),
    .B(_06590_),
    .Y(_06592_)
  );
  NAND _14851_ (
    .A(_01531_),
    .B(_06589_),
    .Y(_06593_)
  );
  NAND _14852_ (
    .A(_06592_),
    .B(_06593_),
    .Y(_06594_)
  );
  OR _14853_ (
    .A(\data_i[0] ),
    .B(_01586_),
    .Y(_06595_)
  );
  AND _14854_ (
    .A(MemWrite_i),
    .B(_06595_),
    .Y(_06596_)
  );
  NAND _14855_ (
    .A(_06594_),
    .B(_06596_),
    .Y(_06597_)
  );
  NAND _14856_ (
    .A(_06583_),
    .B(_06597_),
    .Y(_00216_)
  );
  NAND _14857_ (
    .A(\memory[5][1] ),
    .B(_05361_),
    .Y(_06598_)
  );
  OR _14858_ (
    .A(\memory[5][1] ),
    .B(_01453_),
    .Y(_06599_)
  );
  OR _14859_ (
    .A(\data_i[25] ),
    .B(_01454_),
    .Y(_06600_)
  );
  NAND _14860_ (
    .A(_06599_),
    .B(_06600_),
    .Y(_06602_)
  );
  NAND _14861_ (
    .A(_01514_),
    .B(_06602_),
    .Y(_06603_)
  );
  OR _14862_ (
    .A(\data_i[17] ),
    .B(_01514_),
    .Y(_06604_)
  );
  AND _14863_ (
    .A(_06603_),
    .B(_06604_),
    .Y(_06605_)
  );
  NAND _14864_ (
    .A(\data_i[9] ),
    .B(_01530_),
    .Y(_06606_)
  );
  AND _14865_ (
    .A(_01586_),
    .B(_06606_),
    .Y(_06607_)
  );
  NAND _14866_ (
    .A(_01531_),
    .B(_06605_),
    .Y(_06608_)
  );
  NAND _14867_ (
    .A(_06607_),
    .B(_06608_),
    .Y(_06609_)
  );
  OR _14868_ (
    .A(\data_i[1] ),
    .B(_01586_),
    .Y(_06610_)
  );
  AND _14869_ (
    .A(MemWrite_i),
    .B(_06610_),
    .Y(_06611_)
  );
  NAND _14870_ (
    .A(_06609_),
    .B(_06611_),
    .Y(_06613_)
  );
  NAND _14871_ (
    .A(_06598_),
    .B(_06613_),
    .Y(_00217_)
  );
  NAND _14872_ (
    .A(\memory[5][2] ),
    .B(_05361_),
    .Y(_06614_)
  );
  OR _14873_ (
    .A(\memory[5][2] ),
    .B(_01453_),
    .Y(_06615_)
  );
  OR _14874_ (
    .A(\data_i[26] ),
    .B(_01454_),
    .Y(_06616_)
  );
  NAND _14875_ (
    .A(_06615_),
    .B(_06616_),
    .Y(_06617_)
  );
  NAND _14876_ (
    .A(_01514_),
    .B(_06617_),
    .Y(_06618_)
  );
  OR _14877_ (
    .A(\data_i[18] ),
    .B(_01514_),
    .Y(_06619_)
  );
  AND _14878_ (
    .A(_06618_),
    .B(_06619_),
    .Y(_06620_)
  );
  NAND _14879_ (
    .A(\data_i[10] ),
    .B(_01530_),
    .Y(_06621_)
  );
  AND _14880_ (
    .A(_01586_),
    .B(_06621_),
    .Y(_06623_)
  );
  NAND _14881_ (
    .A(_01531_),
    .B(_06620_),
    .Y(_06624_)
  );
  NAND _14882_ (
    .A(_06623_),
    .B(_06624_),
    .Y(_06625_)
  );
  OR _14883_ (
    .A(\data_i[2] ),
    .B(_01586_),
    .Y(_06626_)
  );
  AND _14884_ (
    .A(MemWrite_i),
    .B(_06626_),
    .Y(_06627_)
  );
  NAND _14885_ (
    .A(_06625_),
    .B(_06627_),
    .Y(_06628_)
  );
  NAND _14886_ (
    .A(_06614_),
    .B(_06628_),
    .Y(_00218_)
  );
  NAND _14887_ (
    .A(\memory[5][3] ),
    .B(_05361_),
    .Y(_06629_)
  );
  OR _14888_ (
    .A(\memory[5][3] ),
    .B(_01453_),
    .Y(_06630_)
  );
  OR _14889_ (
    .A(\data_i[27] ),
    .B(_01454_),
    .Y(_06631_)
  );
  NAND _14890_ (
    .A(_06630_),
    .B(_06631_),
    .Y(_06633_)
  );
  NAND _14891_ (
    .A(_01514_),
    .B(_06633_),
    .Y(_06634_)
  );
  OR _14892_ (
    .A(\data_i[19] ),
    .B(_01514_),
    .Y(_06635_)
  );
  AND _14893_ (
    .A(_06634_),
    .B(_06635_),
    .Y(_06636_)
  );
  NAND _14894_ (
    .A(\data_i[11] ),
    .B(_01530_),
    .Y(_06637_)
  );
  AND _14895_ (
    .A(_01586_),
    .B(_06637_),
    .Y(_06638_)
  );
  NAND _14896_ (
    .A(_01531_),
    .B(_06636_),
    .Y(_06639_)
  );
  NAND _14897_ (
    .A(_06638_),
    .B(_06639_),
    .Y(_06640_)
  );
  OR _14898_ (
    .A(\data_i[3] ),
    .B(_01586_),
    .Y(_06641_)
  );
  AND _14899_ (
    .A(MemWrite_i),
    .B(_06641_),
    .Y(_06642_)
  );
  NAND _14900_ (
    .A(_06640_),
    .B(_06642_),
    .Y(_06644_)
  );
  NAND _14901_ (
    .A(_06629_),
    .B(_06644_),
    .Y(_00219_)
  );
  NAND _14902_ (
    .A(\memory[5][4] ),
    .B(_05361_),
    .Y(_06645_)
  );
  OR _14903_ (
    .A(\memory[5][4] ),
    .B(_01453_),
    .Y(_06646_)
  );
  OR _14904_ (
    .A(\data_i[28] ),
    .B(_01454_),
    .Y(_06647_)
  );
  NAND _14905_ (
    .A(_06646_),
    .B(_06647_),
    .Y(_06648_)
  );
  NAND _14906_ (
    .A(_01514_),
    .B(_06648_),
    .Y(_06649_)
  );
  OR _14907_ (
    .A(\data_i[20] ),
    .B(_01514_),
    .Y(_06650_)
  );
  AND _14908_ (
    .A(_06649_),
    .B(_06650_),
    .Y(_06651_)
  );
  NAND _14909_ (
    .A(\data_i[12] ),
    .B(_01530_),
    .Y(_06652_)
  );
  AND _14910_ (
    .A(_01586_),
    .B(_06652_),
    .Y(_06654_)
  );
  NAND _14911_ (
    .A(_01531_),
    .B(_06651_),
    .Y(_06655_)
  );
  NAND _14912_ (
    .A(_06654_),
    .B(_06655_),
    .Y(_06656_)
  );
  OR _14913_ (
    .A(\data_i[4] ),
    .B(_01586_),
    .Y(_06657_)
  );
  AND _14914_ (
    .A(MemWrite_i),
    .B(_06657_),
    .Y(_06658_)
  );
  NAND _14915_ (
    .A(_06656_),
    .B(_06658_),
    .Y(_06659_)
  );
  NAND _14916_ (
    .A(_06645_),
    .B(_06659_),
    .Y(_00220_)
  );
  NAND _14917_ (
    .A(\memory[5][5] ),
    .B(_05361_),
    .Y(_06660_)
  );
  OR _14918_ (
    .A(\memory[5][5] ),
    .B(_01453_),
    .Y(_06661_)
  );
  OR _14919_ (
    .A(\data_i[29] ),
    .B(_01454_),
    .Y(_06662_)
  );
  NAND _14920_ (
    .A(_06661_),
    .B(_06662_),
    .Y(_06664_)
  );
  NAND _14921_ (
    .A(_01514_),
    .B(_06664_),
    .Y(_06665_)
  );
  OR _14922_ (
    .A(\data_i[21] ),
    .B(_01514_),
    .Y(_06666_)
  );
  AND _14923_ (
    .A(_06665_),
    .B(_06666_),
    .Y(_06667_)
  );
  NAND _14924_ (
    .A(\data_i[13] ),
    .B(_01530_),
    .Y(_06668_)
  );
  AND _14925_ (
    .A(_01586_),
    .B(_06668_),
    .Y(_06669_)
  );
  NAND _14926_ (
    .A(_01531_),
    .B(_06667_),
    .Y(_06670_)
  );
  NAND _14927_ (
    .A(_06669_),
    .B(_06670_),
    .Y(_06671_)
  );
  OR _14928_ (
    .A(\data_i[5] ),
    .B(_01586_),
    .Y(_06672_)
  );
  AND _14929_ (
    .A(MemWrite_i),
    .B(_06672_),
    .Y(_06673_)
  );
  NAND _14930_ (
    .A(_06671_),
    .B(_06673_),
    .Y(_06675_)
  );
  NAND _14931_ (
    .A(_06660_),
    .B(_06675_),
    .Y(_00221_)
  );
  NAND _14932_ (
    .A(\memory[5][6] ),
    .B(_05361_),
    .Y(_06676_)
  );
  OR _14933_ (
    .A(\memory[5][6] ),
    .B(_01453_),
    .Y(_06677_)
  );
  OR _14934_ (
    .A(\data_i[30] ),
    .B(_01454_),
    .Y(_06678_)
  );
  NAND _14935_ (
    .A(_06677_),
    .B(_06678_),
    .Y(_06679_)
  );
  NAND _14936_ (
    .A(_01514_),
    .B(_06679_),
    .Y(_06680_)
  );
  OR _14937_ (
    .A(\data_i[22] ),
    .B(_01514_),
    .Y(_06681_)
  );
  AND _14938_ (
    .A(_06680_),
    .B(_06681_),
    .Y(_06682_)
  );
  NAND _14939_ (
    .A(\data_i[14] ),
    .B(_01530_),
    .Y(_06683_)
  );
  AND _14940_ (
    .A(_01586_),
    .B(_06683_),
    .Y(_06685_)
  );
  NAND _14941_ (
    .A(_01531_),
    .B(_06682_),
    .Y(_06686_)
  );
  NAND _14942_ (
    .A(_06685_),
    .B(_06686_),
    .Y(_06687_)
  );
  OR _14943_ (
    .A(\data_i[6] ),
    .B(_01586_),
    .Y(_06688_)
  );
  AND _14944_ (
    .A(MemWrite_i),
    .B(_06688_),
    .Y(_06689_)
  );
  NAND _14945_ (
    .A(_06687_),
    .B(_06689_),
    .Y(_06690_)
  );
  NAND _14946_ (
    .A(_06676_),
    .B(_06690_),
    .Y(_00222_)
  );
  NAND _14947_ (
    .A(\memory[5][7] ),
    .B(_05361_),
    .Y(_06691_)
  );
  OR _14948_ (
    .A(\memory[5][7] ),
    .B(_01453_),
    .Y(_06692_)
  );
  OR _14949_ (
    .A(\data_i[31] ),
    .B(_01454_),
    .Y(_06693_)
  );
  NAND _14950_ (
    .A(_06692_),
    .B(_06693_),
    .Y(_06695_)
  );
  NAND _14951_ (
    .A(_01514_),
    .B(_06695_),
    .Y(_06696_)
  );
  OR _14952_ (
    .A(\data_i[23] ),
    .B(_01514_),
    .Y(_06697_)
  );
  AND _14953_ (
    .A(_06696_),
    .B(_06697_),
    .Y(_06698_)
  );
  NAND _14954_ (
    .A(\data_i[15] ),
    .B(_01530_),
    .Y(_06699_)
  );
  AND _14955_ (
    .A(_01586_),
    .B(_06699_),
    .Y(_06700_)
  );
  NAND _14956_ (
    .A(_01531_),
    .B(_06698_),
    .Y(_06701_)
  );
  NAND _14957_ (
    .A(_06700_),
    .B(_06701_),
    .Y(_06702_)
  );
  OR _14958_ (
    .A(\data_i[7] ),
    .B(_01586_),
    .Y(_06703_)
  );
  AND _14959_ (
    .A(MemWrite_i),
    .B(_06703_),
    .Y(_06704_)
  );
  NAND _14960_ (
    .A(_06702_),
    .B(_06704_),
    .Y(_06706_)
  );
  NAND _14961_ (
    .A(_06691_),
    .B(_06706_),
    .Y(_00223_)
  );
  OR _14962_ (
    .A(\memory[4][0] ),
    .B(MemWrite_i),
    .Y(_06707_)
  );
  NAND _14963_ (
    .A(\data_i[24] ),
    .B(_01570_),
    .Y(_06708_)
  );
  NAND _14964_ (
    .A(\memory[4][0] ),
    .B(_01571_),
    .Y(_06709_)
  );
  NAND _14965_ (
    .A(_06708_),
    .B(_06709_),
    .Y(_06710_)
  );
  NAND _14966_ (
    .A(_01454_),
    .B(_06710_),
    .Y(_06711_)
  );
  NAND _14967_ (
    .A(\data_i[16] ),
    .B(_01453_),
    .Y(_06712_)
  );
  AND _14968_ (
    .A(_01514_),
    .B(_06712_),
    .Y(_06713_)
  );
  NAND _14969_ (
    .A(_06711_),
    .B(_06713_),
    .Y(_06714_)
  );
  OR _14970_ (
    .A(\data_i[8] ),
    .B(_01514_),
    .Y(_06716_)
  );
  AND _14971_ (
    .A(_01531_),
    .B(_06716_),
    .Y(_06717_)
  );
  NAND _14972_ (
    .A(_06714_),
    .B(_06717_),
    .Y(_06718_)
  );
  NAND _14973_ (
    .A(\data_i[0] ),
    .B(_01530_),
    .Y(_06719_)
  );
  AND _14974_ (
    .A(MemWrite_i),
    .B(_06719_),
    .Y(_06720_)
  );
  NAND _14975_ (
    .A(_06718_),
    .B(_06720_),
    .Y(_06721_)
  );
  AND _14976_ (
    .A(_06707_),
    .B(_06721_),
    .Y(_00208_)
  );
  NAND _14977_ (
    .A(\memory[4][1] ),
    .B(_05361_),
    .Y(_06722_)
  );
  OR _14978_ (
    .A(\memory[4][1] ),
    .B(_01570_),
    .Y(_06723_)
  );
  OR _14979_ (
    .A(\data_i[25] ),
    .B(_01571_),
    .Y(_06724_)
  );
  NAND _14980_ (
    .A(_06723_),
    .B(_06724_),
    .Y(_06725_)
  );
  NAND _14981_ (
    .A(_01454_),
    .B(_06725_),
    .Y(_06726_)
  );
  OR _14982_ (
    .A(\data_i[17] ),
    .B(_01454_),
    .Y(_06727_)
  );
  AND _14983_ (
    .A(_06726_),
    .B(_06727_),
    .Y(_06728_)
  );
  NAND _14984_ (
    .A(\data_i[9] ),
    .B(_01513_),
    .Y(_06729_)
  );
  AND _14985_ (
    .A(_01531_),
    .B(_06729_),
    .Y(_06730_)
  );
  NAND _14986_ (
    .A(_01514_),
    .B(_06728_),
    .Y(_06731_)
  );
  NAND _14987_ (
    .A(_06730_),
    .B(_06731_),
    .Y(_06732_)
  );
  OR _14988_ (
    .A(\data_i[1] ),
    .B(_01531_),
    .Y(_06733_)
  );
  AND _14989_ (
    .A(MemWrite_i),
    .B(_06733_),
    .Y(_06734_)
  );
  NAND _14990_ (
    .A(_06732_),
    .B(_06734_),
    .Y(_06736_)
  );
  NAND _14991_ (
    .A(_06722_),
    .B(_06736_),
    .Y(_00209_)
  );
  NAND _14992_ (
    .A(\memory[4][2] ),
    .B(_05361_),
    .Y(_06737_)
  );
  OR _14993_ (
    .A(\memory[4][2] ),
    .B(_01570_),
    .Y(_06738_)
  );
  OR _14994_ (
    .A(\data_i[26] ),
    .B(_01571_),
    .Y(_06739_)
  );
  NAND _14995_ (
    .A(_06738_),
    .B(_06739_),
    .Y(_06740_)
  );
  NAND _14996_ (
    .A(_01454_),
    .B(_06740_),
    .Y(_06741_)
  );
  OR _14997_ (
    .A(\data_i[18] ),
    .B(_01454_),
    .Y(_06742_)
  );
  AND _14998_ (
    .A(_06741_),
    .B(_06742_),
    .Y(_06743_)
  );
  NAND _14999_ (
    .A(\data_i[10] ),
    .B(_01513_),
    .Y(_06744_)
  );
  AND _15000_ (
    .A(_01531_),
    .B(_06744_),
    .Y(_06746_)
  );
  NAND _15001_ (
    .A(_01514_),
    .B(_06743_),
    .Y(_06747_)
  );
  NAND _15002_ (
    .A(_06746_),
    .B(_06747_),
    .Y(_06748_)
  );
  OR _15003_ (
    .A(\data_i[2] ),
    .B(_01531_),
    .Y(_06749_)
  );
  AND _15004_ (
    .A(MemWrite_i),
    .B(_06749_),
    .Y(_06750_)
  );
  NAND _15005_ (
    .A(_06748_),
    .B(_06750_),
    .Y(_06751_)
  );
  NAND _15006_ (
    .A(_06737_),
    .B(_06751_),
    .Y(_00210_)
  );
  NAND _15007_ (
    .A(\memory[4][3] ),
    .B(_05361_),
    .Y(_06752_)
  );
  OR _15008_ (
    .A(\memory[4][3] ),
    .B(_01570_),
    .Y(_06753_)
  );
  OR _15009_ (
    .A(\data_i[27] ),
    .B(_01571_),
    .Y(_06754_)
  );
  NAND _15010_ (
    .A(_06753_),
    .B(_06754_),
    .Y(_06756_)
  );
  NAND _15011_ (
    .A(_01454_),
    .B(_06756_),
    .Y(_06757_)
  );
  OR _15012_ (
    .A(\data_i[19] ),
    .B(_01454_),
    .Y(_06758_)
  );
  AND _15013_ (
    .A(_06757_),
    .B(_06758_),
    .Y(_06759_)
  );
  NAND _15014_ (
    .A(\data_i[11] ),
    .B(_01513_),
    .Y(_06760_)
  );
  AND _15015_ (
    .A(_01531_),
    .B(_06760_),
    .Y(_06761_)
  );
  NAND _15016_ (
    .A(_01514_),
    .B(_06759_),
    .Y(_06762_)
  );
  NAND _15017_ (
    .A(_06761_),
    .B(_06762_),
    .Y(_06763_)
  );
  OR _15018_ (
    .A(\data_i[3] ),
    .B(_01531_),
    .Y(_06764_)
  );
  AND _15019_ (
    .A(MemWrite_i),
    .B(_06764_),
    .Y(_06765_)
  );
  NAND _15020_ (
    .A(_06763_),
    .B(_06765_),
    .Y(_06767_)
  );
  NAND _15021_ (
    .A(_06752_),
    .B(_06767_),
    .Y(_00211_)
  );
  NAND _15022_ (
    .A(\memory[4][4] ),
    .B(_05361_),
    .Y(_06768_)
  );
  OR _15023_ (
    .A(\memory[4][4] ),
    .B(_01570_),
    .Y(_06769_)
  );
  OR _15024_ (
    .A(\data_i[28] ),
    .B(_01571_),
    .Y(_06770_)
  );
  NAND _15025_ (
    .A(_06769_),
    .B(_06770_),
    .Y(_06771_)
  );
  NAND _15026_ (
    .A(_01454_),
    .B(_06771_),
    .Y(_06772_)
  );
  OR _15027_ (
    .A(\data_i[20] ),
    .B(_01454_),
    .Y(_06773_)
  );
  AND _15028_ (
    .A(_06772_),
    .B(_06773_),
    .Y(_06774_)
  );
  NAND _15029_ (
    .A(\data_i[12] ),
    .B(_01513_),
    .Y(_06775_)
  );
  AND _15030_ (
    .A(_01531_),
    .B(_06775_),
    .Y(_06777_)
  );
  NAND _15031_ (
    .A(_01514_),
    .B(_06774_),
    .Y(_06778_)
  );
  NAND _15032_ (
    .A(_06777_),
    .B(_06778_),
    .Y(_06779_)
  );
  OR _15033_ (
    .A(\data_i[4] ),
    .B(_01531_),
    .Y(_06780_)
  );
  AND _15034_ (
    .A(MemWrite_i),
    .B(_06780_),
    .Y(_06781_)
  );
  NAND _15035_ (
    .A(_06779_),
    .B(_06781_),
    .Y(_06782_)
  );
  NAND _15036_ (
    .A(_06768_),
    .B(_06782_),
    .Y(_00212_)
  );
  NAND _15037_ (
    .A(\memory[4][5] ),
    .B(_05361_),
    .Y(_06783_)
  );
  OR _15038_ (
    .A(\memory[4][5] ),
    .B(_01570_),
    .Y(_06784_)
  );
  OR _15039_ (
    .A(\data_i[29] ),
    .B(_01571_),
    .Y(_06785_)
  );
  NAND _15040_ (
    .A(_06784_),
    .B(_06785_),
    .Y(_06787_)
  );
  NAND _15041_ (
    .A(_01454_),
    .B(_06787_),
    .Y(_06788_)
  );
  OR _15042_ (
    .A(\data_i[21] ),
    .B(_01454_),
    .Y(_06789_)
  );
  AND _15043_ (
    .A(_06788_),
    .B(_06789_),
    .Y(_06790_)
  );
  NAND _15044_ (
    .A(\data_i[13] ),
    .B(_01513_),
    .Y(_06791_)
  );
  AND _15045_ (
    .A(_01531_),
    .B(_06791_),
    .Y(_06792_)
  );
  NAND _15046_ (
    .A(_01514_),
    .B(_06790_),
    .Y(_06793_)
  );
  NAND _15047_ (
    .A(_06792_),
    .B(_06793_),
    .Y(_06794_)
  );
  OR _15048_ (
    .A(\data_i[5] ),
    .B(_01531_),
    .Y(_06795_)
  );
  AND _15049_ (
    .A(MemWrite_i),
    .B(_06795_),
    .Y(_06796_)
  );
  NAND _15050_ (
    .A(_06794_),
    .B(_06796_),
    .Y(_06798_)
  );
  NAND _15051_ (
    .A(_06783_),
    .B(_06798_),
    .Y(_00213_)
  );
  NAND _15052_ (
    .A(\memory[4][6] ),
    .B(_05361_),
    .Y(_06799_)
  );
  OR _15053_ (
    .A(\memory[4][6] ),
    .B(_01570_),
    .Y(_06800_)
  );
  OR _15054_ (
    .A(\data_i[30] ),
    .B(_01571_),
    .Y(_06801_)
  );
  NAND _15055_ (
    .A(_06800_),
    .B(_06801_),
    .Y(_06802_)
  );
  NAND _15056_ (
    .A(_01454_),
    .B(_06802_),
    .Y(_06803_)
  );
  OR _15057_ (
    .A(\data_i[22] ),
    .B(_01454_),
    .Y(_06804_)
  );
  AND _15058_ (
    .A(_06803_),
    .B(_06804_),
    .Y(_06805_)
  );
  NAND _15059_ (
    .A(\data_i[14] ),
    .B(_01513_),
    .Y(_06806_)
  );
  AND _15060_ (
    .A(_01531_),
    .B(_06806_),
    .Y(_06808_)
  );
  NAND _15061_ (
    .A(_01514_),
    .B(_06805_),
    .Y(_06809_)
  );
  NAND _15062_ (
    .A(_06808_),
    .B(_06809_),
    .Y(_06810_)
  );
  OR _15063_ (
    .A(\data_i[6] ),
    .B(_01531_),
    .Y(_06811_)
  );
  AND _15064_ (
    .A(MemWrite_i),
    .B(_06811_),
    .Y(_06812_)
  );
  NAND _15065_ (
    .A(_06810_),
    .B(_06812_),
    .Y(_06813_)
  );
  NAND _15066_ (
    .A(_06799_),
    .B(_06813_),
    .Y(_00214_)
  );
  NAND _15067_ (
    .A(\memory[4][7] ),
    .B(_05361_),
    .Y(_06814_)
  );
  OR _15068_ (
    .A(\memory[4][7] ),
    .B(_01570_),
    .Y(_06815_)
  );
  OR _15069_ (
    .A(\data_i[31] ),
    .B(_01571_),
    .Y(_06816_)
  );
  NAND _15070_ (
    .A(_06815_),
    .B(_06816_),
    .Y(_06818_)
  );
  NAND _15071_ (
    .A(_01454_),
    .B(_06818_),
    .Y(_06819_)
  );
  OR _15072_ (
    .A(\data_i[23] ),
    .B(_01454_),
    .Y(_06820_)
  );
  AND _15073_ (
    .A(_06819_),
    .B(_06820_),
    .Y(_06821_)
  );
  NAND _15074_ (
    .A(\data_i[15] ),
    .B(_01513_),
    .Y(_06822_)
  );
  AND _15075_ (
    .A(_01531_),
    .B(_06822_),
    .Y(_06823_)
  );
  NAND _15076_ (
    .A(_01514_),
    .B(_06821_),
    .Y(_06824_)
  );
  NAND _15077_ (
    .A(_06823_),
    .B(_06824_),
    .Y(_06825_)
  );
  OR _15078_ (
    .A(\data_i[7] ),
    .B(_01531_),
    .Y(_06826_)
  );
  AND _15079_ (
    .A(MemWrite_i),
    .B(_06826_),
    .Y(_06827_)
  );
  NAND _15080_ (
    .A(_06825_),
    .B(_06827_),
    .Y(_06829_)
  );
  NAND _15081_ (
    .A(_06814_),
    .B(_06829_),
    .Y(_00215_)
  );
  NAND _15082_ (
    .A(\memory[3][0] ),
    .B(_05361_),
    .Y(_06830_)
  );
  OR _15083_ (
    .A(\memory[3][0] ),
    .B(_01449_),
    .Y(_06831_)
  );
  OR _15084_ (
    .A(\data_i[24] ),
    .B(_01450_),
    .Y(_06832_)
  );
  NAND _15085_ (
    .A(_06831_),
    .B(_06832_),
    .Y(_06833_)
  );
  NAND _15086_ (
    .A(_01571_),
    .B(_06833_),
    .Y(_06834_)
  );
  OR _15087_ (
    .A(\data_i[16] ),
    .B(_01571_),
    .Y(_06835_)
  );
  AND _15088_ (
    .A(_06834_),
    .B(_06835_),
    .Y(_06836_)
  );
  NAND _15089_ (
    .A(\data_i[8] ),
    .B(_01453_),
    .Y(_06837_)
  );
  AND _15090_ (
    .A(_01514_),
    .B(_06837_),
    .Y(_06839_)
  );
  NAND _15091_ (
    .A(_01454_),
    .B(_06836_),
    .Y(_06840_)
  );
  NAND _15092_ (
    .A(_06839_),
    .B(_06840_),
    .Y(_06841_)
  );
  OR _15093_ (
    .A(\data_i[0] ),
    .B(_01514_),
    .Y(_06842_)
  );
  AND _15094_ (
    .A(MemWrite_i),
    .B(_06842_),
    .Y(_06843_)
  );
  NAND _15095_ (
    .A(_06841_),
    .B(_06843_),
    .Y(_06844_)
  );
  NAND _15096_ (
    .A(_06830_),
    .B(_06844_),
    .Y(_00200_)
  );
  OR _15097_ (
    .A(\memory[3][1] ),
    .B(MemWrite_i),
    .Y(_06845_)
  );
  NAND _15098_ (
    .A(\data_i[25] ),
    .B(_01449_),
    .Y(_06846_)
  );
  NAND _15099_ (
    .A(\memory[3][1] ),
    .B(_01450_),
    .Y(_06847_)
  );
  NAND _15100_ (
    .A(_06846_),
    .B(_06847_),
    .Y(_06849_)
  );
  NAND _15101_ (
    .A(_01571_),
    .B(_06849_),
    .Y(_06850_)
  );
  NAND _15102_ (
    .A(\data_i[17] ),
    .B(_01570_),
    .Y(_06851_)
  );
  AND _15103_ (
    .A(_06850_),
    .B(_06851_),
    .Y(_06852_)
  );
  OR _15104_ (
    .A(\data_i[9] ),
    .B(_01454_),
    .Y(_06853_)
  );
  AND _15105_ (
    .A(_01514_),
    .B(_06853_),
    .Y(_06854_)
  );
  NAND _15106_ (
    .A(_01454_),
    .B(_06852_),
    .Y(_06855_)
  );
  NAND _15107_ (
    .A(_06854_),
    .B(_06855_),
    .Y(_06856_)
  );
  NAND _15108_ (
    .A(\data_i[1] ),
    .B(_01513_),
    .Y(_06857_)
  );
  AND _15109_ (
    .A(MemWrite_i),
    .B(_06857_),
    .Y(_06858_)
  );
  NAND _15110_ (
    .A(_06856_),
    .B(_06858_),
    .Y(_06860_)
  );
  AND _15111_ (
    .A(_06845_),
    .B(_06860_),
    .Y(_00201_)
  );
  OR _15112_ (
    .A(\memory[3][2] ),
    .B(MemWrite_i),
    .Y(_06861_)
  );
  NAND _15113_ (
    .A(\data_i[26] ),
    .B(_01449_),
    .Y(_06862_)
  );
  NAND _15114_ (
    .A(\memory[3][2] ),
    .B(_01450_),
    .Y(_06863_)
  );
  NAND _15115_ (
    .A(_06862_),
    .B(_06863_),
    .Y(_06864_)
  );
  NAND _15116_ (
    .A(_01571_),
    .B(_06864_),
    .Y(_06865_)
  );
  NAND _15117_ (
    .A(\data_i[18] ),
    .B(_01570_),
    .Y(_06866_)
  );
  AND _15118_ (
    .A(_01454_),
    .B(_06866_),
    .Y(_06867_)
  );
  NAND _15119_ (
    .A(_06865_),
    .B(_06867_),
    .Y(_06868_)
  );
  OR _15120_ (
    .A(\data_i[10] ),
    .B(_01454_),
    .Y(_06870_)
  );
  AND _15121_ (
    .A(_01514_),
    .B(_06870_),
    .Y(_06871_)
  );
  NAND _15122_ (
    .A(_06868_),
    .B(_06871_),
    .Y(_06872_)
  );
  NAND _15123_ (
    .A(\data_i[2] ),
    .B(_01513_),
    .Y(_06873_)
  );
  AND _15124_ (
    .A(MemWrite_i),
    .B(_06873_),
    .Y(_06874_)
  );
  NAND _15125_ (
    .A(_06872_),
    .B(_06874_),
    .Y(_06875_)
  );
  AND _15126_ (
    .A(_06861_),
    .B(_06875_),
    .Y(_00202_)
  );
  NAND _15127_ (
    .A(\memory[3][3] ),
    .B(_05361_),
    .Y(_06876_)
  );
  OR _15128_ (
    .A(\memory[3][3] ),
    .B(_01449_),
    .Y(_06877_)
  );
  OR _15129_ (
    .A(\data_i[27] ),
    .B(_01450_),
    .Y(_06878_)
  );
  NAND _15130_ (
    .A(_06877_),
    .B(_06878_),
    .Y(_06880_)
  );
  NAND _15131_ (
    .A(_01571_),
    .B(_06880_),
    .Y(_06881_)
  );
  OR _15132_ (
    .A(\data_i[19] ),
    .B(_01571_),
    .Y(_06882_)
  );
  AND _15133_ (
    .A(_06881_),
    .B(_06882_),
    .Y(_06883_)
  );
  NAND _15134_ (
    .A(\data_i[11] ),
    .B(_01453_),
    .Y(_06884_)
  );
  AND _15135_ (
    .A(_01514_),
    .B(_06884_),
    .Y(_06885_)
  );
  NAND _15136_ (
    .A(_01454_),
    .B(_06883_),
    .Y(_06886_)
  );
  NAND _15137_ (
    .A(_06885_),
    .B(_06886_),
    .Y(_06887_)
  );
  OR _15138_ (
    .A(\data_i[3] ),
    .B(_01514_),
    .Y(_06888_)
  );
  AND _15139_ (
    .A(MemWrite_i),
    .B(_06888_),
    .Y(_06889_)
  );
  NAND _15140_ (
    .A(_06887_),
    .B(_06889_),
    .Y(_06891_)
  );
  NAND _15141_ (
    .A(_06876_),
    .B(_06891_),
    .Y(_00203_)
  );
  OR _15142_ (
    .A(\memory[3][4] ),
    .B(MemWrite_i),
    .Y(_06892_)
  );
  NAND _15143_ (
    .A(\data_i[28] ),
    .B(_01449_),
    .Y(_06893_)
  );
  NAND _15144_ (
    .A(\memory[3][4] ),
    .B(_01450_),
    .Y(_06894_)
  );
  NAND _15145_ (
    .A(_06893_),
    .B(_06894_),
    .Y(_06895_)
  );
  NAND _15146_ (
    .A(_01571_),
    .B(_06895_),
    .Y(_06896_)
  );
  NAND _15147_ (
    .A(\data_i[20] ),
    .B(_01570_),
    .Y(_06897_)
  );
  AND _15148_ (
    .A(_01454_),
    .B(_06897_),
    .Y(_06898_)
  );
  NAND _15149_ (
    .A(_06896_),
    .B(_06898_),
    .Y(_06899_)
  );
  OR _15150_ (
    .A(\data_i[12] ),
    .B(_01454_),
    .Y(_06901_)
  );
  AND _15151_ (
    .A(_01514_),
    .B(_06901_),
    .Y(_06902_)
  );
  NAND _15152_ (
    .A(_06899_),
    .B(_06902_),
    .Y(_06903_)
  );
  NAND _15153_ (
    .A(\data_i[4] ),
    .B(_01513_),
    .Y(_06904_)
  );
  AND _15154_ (
    .A(MemWrite_i),
    .B(_06904_),
    .Y(_06905_)
  );
  NAND _15155_ (
    .A(_06903_),
    .B(_06905_),
    .Y(_06906_)
  );
  AND _15156_ (
    .A(_06892_),
    .B(_06906_),
    .Y(_00204_)
  );
  NAND _15157_ (
    .A(\memory[3][5] ),
    .B(_05361_),
    .Y(_06907_)
  );
  OR _15158_ (
    .A(\memory[3][5] ),
    .B(_01449_),
    .Y(_06908_)
  );
  OR _15159_ (
    .A(\data_i[29] ),
    .B(_01450_),
    .Y(_06909_)
  );
  NAND _15160_ (
    .A(_06908_),
    .B(_06909_),
    .Y(_06911_)
  );
  NAND _15161_ (
    .A(_01571_),
    .B(_06911_),
    .Y(_06912_)
  );
  OR _15162_ (
    .A(\data_i[21] ),
    .B(_01571_),
    .Y(_06913_)
  );
  AND _15163_ (
    .A(_06912_),
    .B(_06913_),
    .Y(_06914_)
  );
  NAND _15164_ (
    .A(\data_i[13] ),
    .B(_01453_),
    .Y(_06915_)
  );
  AND _15165_ (
    .A(_01514_),
    .B(_06915_),
    .Y(_06916_)
  );
  NAND _15166_ (
    .A(_01454_),
    .B(_06914_),
    .Y(_06917_)
  );
  NAND _15167_ (
    .A(_06916_),
    .B(_06917_),
    .Y(_06918_)
  );
  OR _15168_ (
    .A(\data_i[5] ),
    .B(_01514_),
    .Y(_06919_)
  );
  AND _15169_ (
    .A(MemWrite_i),
    .B(_06919_),
    .Y(_06920_)
  );
  NAND _15170_ (
    .A(_06918_),
    .B(_06920_),
    .Y(_06922_)
  );
  NAND _15171_ (
    .A(_06907_),
    .B(_06922_),
    .Y(_00205_)
  );
  NAND _15172_ (
    .A(\memory[3][6] ),
    .B(_05361_),
    .Y(_06923_)
  );
  OR _15173_ (
    .A(\memory[3][6] ),
    .B(_01449_),
    .Y(_06924_)
  );
  OR _15174_ (
    .A(\data_i[30] ),
    .B(_01450_),
    .Y(_06925_)
  );
  NAND _15175_ (
    .A(_06924_),
    .B(_06925_),
    .Y(_06926_)
  );
  NAND _15176_ (
    .A(_01571_),
    .B(_06926_),
    .Y(_06927_)
  );
  OR _15177_ (
    .A(\data_i[22] ),
    .B(_01571_),
    .Y(_06928_)
  );
  AND _15178_ (
    .A(_06927_),
    .B(_06928_),
    .Y(_06929_)
  );
  NAND _15179_ (
    .A(\data_i[14] ),
    .B(_01453_),
    .Y(_06930_)
  );
  AND _15180_ (
    .A(_01514_),
    .B(_06930_),
    .Y(_06932_)
  );
  NAND _15181_ (
    .A(_01454_),
    .B(_06929_),
    .Y(_06933_)
  );
  NAND _15182_ (
    .A(_06932_),
    .B(_06933_),
    .Y(_06934_)
  );
  OR _15183_ (
    .A(\data_i[6] ),
    .B(_01514_),
    .Y(_06935_)
  );
  AND _15184_ (
    .A(MemWrite_i),
    .B(_06935_),
    .Y(_06936_)
  );
  NAND _15185_ (
    .A(_06934_),
    .B(_06936_),
    .Y(_06937_)
  );
  NAND _15186_ (
    .A(_06923_),
    .B(_06937_),
    .Y(_00206_)
  );
  NAND _15187_ (
    .A(\memory[3][7] ),
    .B(_05361_),
    .Y(_06938_)
  );
  OR _15188_ (
    .A(\memory[3][7] ),
    .B(_01449_),
    .Y(_06939_)
  );
  OR _15189_ (
    .A(\data_i[31] ),
    .B(_01450_),
    .Y(_06940_)
  );
  NAND _15190_ (
    .A(_06939_),
    .B(_06940_),
    .Y(_06942_)
  );
  NAND _15191_ (
    .A(_01571_),
    .B(_06942_),
    .Y(_06943_)
  );
  OR _15192_ (
    .A(\data_i[23] ),
    .B(_01571_),
    .Y(_06944_)
  );
  AND _15193_ (
    .A(_06943_),
    .B(_06944_),
    .Y(_06945_)
  );
  NAND _15194_ (
    .A(\data_i[15] ),
    .B(_01453_),
    .Y(_06946_)
  );
  AND _15195_ (
    .A(_01514_),
    .B(_06946_),
    .Y(_06947_)
  );
  NAND _15196_ (
    .A(_01454_),
    .B(_06945_),
    .Y(_06948_)
  );
  NAND _15197_ (
    .A(_06947_),
    .B(_06948_),
    .Y(_06949_)
  );
  OR _15198_ (
    .A(\data_i[7] ),
    .B(_01514_),
    .Y(_06950_)
  );
  AND _15199_ (
    .A(MemWrite_i),
    .B(_06950_),
    .Y(_06951_)
  );
  NAND _15200_ (
    .A(_06949_),
    .B(_06951_),
    .Y(_06953_)
  );
  NAND _15201_ (
    .A(_06938_),
    .B(_06953_),
    .Y(_00207_)
  );
  OR _15202_ (
    .A(\memory[2][0] ),
    .B(MemWrite_i),
    .Y(_06954_)
  );
  NAND _15203_ (
    .A(\data_i[24] ),
    .B(_01504_),
    .Y(_06955_)
  );
  NAND _15204_ (
    .A(\memory[2][0] ),
    .B(_01505_),
    .Y(_06956_)
  );
  NAND _15205_ (
    .A(_06955_),
    .B(_06956_),
    .Y(_06957_)
  );
  NAND _15206_ (
    .A(_01450_),
    .B(_06957_),
    .Y(_06958_)
  );
  NAND _15207_ (
    .A(\data_i[16] ),
    .B(_01449_),
    .Y(_06959_)
  );
  AND _15208_ (
    .A(_01571_),
    .B(_06959_),
    .Y(_06960_)
  );
  NAND _15209_ (
    .A(_06958_),
    .B(_06960_),
    .Y(_06961_)
  );
  OR _15210_ (
    .A(\data_i[8] ),
    .B(_01571_),
    .Y(_06963_)
  );
  AND _15211_ (
    .A(_01454_),
    .B(_06963_),
    .Y(_06964_)
  );
  NAND _15212_ (
    .A(_06961_),
    .B(_06964_),
    .Y(_06965_)
  );
  NAND _15213_ (
    .A(\data_i[0] ),
    .B(_01453_),
    .Y(_06966_)
  );
  AND _15214_ (
    .A(MemWrite_i),
    .B(_06966_),
    .Y(_06967_)
  );
  NAND _15215_ (
    .A(_06965_),
    .B(_06967_),
    .Y(_06968_)
  );
  AND _15216_ (
    .A(_06954_),
    .B(_06968_),
    .Y(_00176_)
  );
  OR _15217_ (
    .A(\memory[2][1] ),
    .B(MemWrite_i),
    .Y(_06969_)
  );
  NAND _15218_ (
    .A(\data_i[25] ),
    .B(_01504_),
    .Y(_06970_)
  );
  NAND _15219_ (
    .A(\memory[2][1] ),
    .B(_01505_),
    .Y(_06971_)
  );
  NAND _15220_ (
    .A(_06970_),
    .B(_06971_),
    .Y(_06973_)
  );
  NAND _15221_ (
    .A(_01450_),
    .B(_06973_),
    .Y(_06974_)
  );
  NAND _15222_ (
    .A(\data_i[17] ),
    .B(_01449_),
    .Y(_06975_)
  );
  AND _15223_ (
    .A(_01571_),
    .B(_06975_),
    .Y(_06976_)
  );
  NAND _15224_ (
    .A(_06974_),
    .B(_06976_),
    .Y(_06977_)
  );
  OR _15225_ (
    .A(\data_i[9] ),
    .B(_01571_),
    .Y(_06978_)
  );
  AND _15226_ (
    .A(_01454_),
    .B(_06978_),
    .Y(_06979_)
  );
  NAND _15227_ (
    .A(_06977_),
    .B(_06979_),
    .Y(_06980_)
  );
  NAND _15228_ (
    .A(\data_i[1] ),
    .B(_01453_),
    .Y(_06981_)
  );
  AND _15229_ (
    .A(MemWrite_i),
    .B(_06981_),
    .Y(_06982_)
  );
  NAND _15230_ (
    .A(_06980_),
    .B(_06982_),
    .Y(_06984_)
  );
  AND _15231_ (
    .A(_06969_),
    .B(_06984_),
    .Y(_00177_)
  );
  NAND _15232_ (
    .A(\memory[2][2] ),
    .B(_05361_),
    .Y(_06985_)
  );
  OR _15233_ (
    .A(\memory[2][2] ),
    .B(_01504_),
    .Y(_06986_)
  );
  OR _15234_ (
    .A(\data_i[26] ),
    .B(_01505_),
    .Y(_06987_)
  );
  NAND _15235_ (
    .A(_06986_),
    .B(_06987_),
    .Y(_06988_)
  );
  NAND _15236_ (
    .A(_01450_),
    .B(_06988_),
    .Y(_06989_)
  );
  OR _15237_ (
    .A(\data_i[18] ),
    .B(_01450_),
    .Y(_06990_)
  );
  AND _15238_ (
    .A(_06989_),
    .B(_06990_),
    .Y(_06991_)
  );
  NAND _15239_ (
    .A(\data_i[10] ),
    .B(_01570_),
    .Y(_06992_)
  );
  AND _15240_ (
    .A(_01454_),
    .B(_06992_),
    .Y(_06994_)
  );
  NAND _15241_ (
    .A(_01571_),
    .B(_06991_),
    .Y(_06995_)
  );
  NAND _15242_ (
    .A(_06994_),
    .B(_06995_),
    .Y(_06996_)
  );
  OR _15243_ (
    .A(\data_i[2] ),
    .B(_01454_),
    .Y(_06997_)
  );
  AND _15244_ (
    .A(MemWrite_i),
    .B(_06997_),
    .Y(_06998_)
  );
  NAND _15245_ (
    .A(_06996_),
    .B(_06998_),
    .Y(_06999_)
  );
  NAND _15246_ (
    .A(_06985_),
    .B(_06999_),
    .Y(_00178_)
  );
  NAND _15247_ (
    .A(\memory[2][3] ),
    .B(_05361_),
    .Y(_07000_)
  );
  OR _15248_ (
    .A(\memory[2][3] ),
    .B(_01504_),
    .Y(_07001_)
  );
  OR _15249_ (
    .A(\data_i[27] ),
    .B(_01505_),
    .Y(_07002_)
  );
  NAND _15250_ (
    .A(_07001_),
    .B(_07002_),
    .Y(_07004_)
  );
  NAND _15251_ (
    .A(_01450_),
    .B(_07004_),
    .Y(_07005_)
  );
  OR _15252_ (
    .A(\data_i[19] ),
    .B(_01450_),
    .Y(_07006_)
  );
  AND _15253_ (
    .A(_07005_),
    .B(_07006_),
    .Y(_07007_)
  );
  NAND _15254_ (
    .A(\data_i[11] ),
    .B(_01570_),
    .Y(_07008_)
  );
  AND _15255_ (
    .A(_01454_),
    .B(_07008_),
    .Y(_07009_)
  );
  NAND _15256_ (
    .A(_01571_),
    .B(_07007_),
    .Y(_07010_)
  );
  NAND _15257_ (
    .A(_07009_),
    .B(_07010_),
    .Y(_07011_)
  );
  OR _15258_ (
    .A(\data_i[3] ),
    .B(_01454_),
    .Y(_07012_)
  );
  AND _15259_ (
    .A(MemWrite_i),
    .B(_07012_),
    .Y(_07013_)
  );
  NAND _15260_ (
    .A(_07011_),
    .B(_07013_),
    .Y(_07015_)
  );
  NAND _15261_ (
    .A(_07000_),
    .B(_07015_),
    .Y(_00179_)
  );
  NAND _15262_ (
    .A(\memory[2][4] ),
    .B(_05361_),
    .Y(_07016_)
  );
  OR _15263_ (
    .A(\memory[2][4] ),
    .B(_01504_),
    .Y(_07017_)
  );
  OR _15264_ (
    .A(\data_i[28] ),
    .B(_01505_),
    .Y(_07018_)
  );
  NAND _15265_ (
    .A(_07017_),
    .B(_07018_),
    .Y(_07019_)
  );
  NAND _15266_ (
    .A(_01450_),
    .B(_07019_),
    .Y(_07020_)
  );
  OR _15267_ (
    .A(\data_i[20] ),
    .B(_01450_),
    .Y(_07021_)
  );
  AND _15268_ (
    .A(_07020_),
    .B(_07021_),
    .Y(_07022_)
  );
  NAND _15269_ (
    .A(\data_i[12] ),
    .B(_01570_),
    .Y(_07023_)
  );
  AND _15270_ (
    .A(_01454_),
    .B(_07023_),
    .Y(_07025_)
  );
  NAND _15271_ (
    .A(_01571_),
    .B(_07022_),
    .Y(_07026_)
  );
  NAND _15272_ (
    .A(_07025_),
    .B(_07026_),
    .Y(_07027_)
  );
  OR _15273_ (
    .A(\data_i[4] ),
    .B(_01454_),
    .Y(_07028_)
  );
  AND _15274_ (
    .A(MemWrite_i),
    .B(_07028_),
    .Y(_07029_)
  );
  NAND _15275_ (
    .A(_07027_),
    .B(_07029_),
    .Y(_07030_)
  );
  NAND _15276_ (
    .A(_07016_),
    .B(_07030_),
    .Y(_00180_)
  );
  NAND _15277_ (
    .A(\memory[2][5] ),
    .B(_05361_),
    .Y(_07031_)
  );
  OR _15278_ (
    .A(\memory[2][5] ),
    .B(_01504_),
    .Y(_07032_)
  );
  OR _15279_ (
    .A(\data_i[29] ),
    .B(_01505_),
    .Y(_07033_)
  );
  NAND _15280_ (
    .A(_07032_),
    .B(_07033_),
    .Y(_07035_)
  );
  NAND _15281_ (
    .A(_01450_),
    .B(_07035_),
    .Y(_07036_)
  );
  OR _15282_ (
    .A(\data_i[21] ),
    .B(_01450_),
    .Y(_07037_)
  );
  AND _15283_ (
    .A(_07036_),
    .B(_07037_),
    .Y(_07038_)
  );
  NAND _15284_ (
    .A(\data_i[13] ),
    .B(_01570_),
    .Y(_07039_)
  );
  AND _15285_ (
    .A(_01454_),
    .B(_07039_),
    .Y(_07040_)
  );
  NAND _15286_ (
    .A(_01571_),
    .B(_07038_),
    .Y(_07041_)
  );
  NAND _15287_ (
    .A(_07040_),
    .B(_07041_),
    .Y(_07042_)
  );
  OR _15288_ (
    .A(\data_i[5] ),
    .B(_01454_),
    .Y(_07043_)
  );
  AND _15289_ (
    .A(MemWrite_i),
    .B(_07043_),
    .Y(_07044_)
  );
  NAND _15290_ (
    .A(_07042_),
    .B(_07044_),
    .Y(_07046_)
  );
  NAND _15291_ (
    .A(_07031_),
    .B(_07046_),
    .Y(_00181_)
  );
  NAND _15292_ (
    .A(\memory[2][6] ),
    .B(_05361_),
    .Y(_07047_)
  );
  OR _15293_ (
    .A(\memory[2][6] ),
    .B(_01504_),
    .Y(_07048_)
  );
  OR _15294_ (
    .A(\data_i[30] ),
    .B(_01505_),
    .Y(_07049_)
  );
  NAND _15295_ (
    .A(_07048_),
    .B(_07049_),
    .Y(_07050_)
  );
  NAND _15296_ (
    .A(_01450_),
    .B(_07050_),
    .Y(_07051_)
  );
  OR _15297_ (
    .A(\data_i[22] ),
    .B(_01450_),
    .Y(_07052_)
  );
  AND _15298_ (
    .A(_07051_),
    .B(_07052_),
    .Y(_07053_)
  );
  NAND _15299_ (
    .A(\data_i[14] ),
    .B(_01570_),
    .Y(_07054_)
  );
  AND _15300_ (
    .A(_01454_),
    .B(_07054_),
    .Y(_07056_)
  );
  NAND _15301_ (
    .A(_01571_),
    .B(_07053_),
    .Y(_07057_)
  );
  NAND _15302_ (
    .A(_07056_),
    .B(_07057_),
    .Y(_07058_)
  );
  OR _15303_ (
    .A(\data_i[6] ),
    .B(_01454_),
    .Y(_07059_)
  );
  AND _15304_ (
    .A(MemWrite_i),
    .B(_07059_),
    .Y(_07060_)
  );
  NAND _15305_ (
    .A(_07058_),
    .B(_07060_),
    .Y(_07061_)
  );
  NAND _15306_ (
    .A(_07047_),
    .B(_07061_),
    .Y(_00182_)
  );
  OR _15307_ (
    .A(\memory[2][7] ),
    .B(MemWrite_i),
    .Y(_07062_)
  );
  NAND _15308_ (
    .A(\data_i[31] ),
    .B(_01504_),
    .Y(_07063_)
  );
  NAND _15309_ (
    .A(\memory[2][7] ),
    .B(_01505_),
    .Y(_07064_)
  );
  NAND _15310_ (
    .A(_07063_),
    .B(_07064_),
    .Y(_07066_)
  );
  NAND _15311_ (
    .A(_01450_),
    .B(_07066_),
    .Y(_07067_)
  );
  NAND _15312_ (
    .A(\data_i[23] ),
    .B(_01449_),
    .Y(_07068_)
  );
  AND _15313_ (
    .A(_07067_),
    .B(_07068_),
    .Y(_07069_)
  );
  OR _15314_ (
    .A(\data_i[15] ),
    .B(_01571_),
    .Y(_07070_)
  );
  AND _15315_ (
    .A(_01454_),
    .B(_07070_),
    .Y(_07071_)
  );
  NAND _15316_ (
    .A(_01571_),
    .B(_07069_),
    .Y(_07072_)
  );
  NAND _15317_ (
    .A(_07071_),
    .B(_07072_),
    .Y(_07073_)
  );
  NAND _15318_ (
    .A(\data_i[7] ),
    .B(_01453_),
    .Y(_07074_)
  );
  AND _15319_ (
    .A(MemWrite_i),
    .B(_07074_),
    .Y(_07075_)
  );
  NAND _15320_ (
    .A(_07073_),
    .B(_07075_),
    .Y(_07077_)
  );
  AND _15321_ (
    .A(_07062_),
    .B(_07077_),
    .Y(_00183_)
  );
  NAND _15322_ (
    .A(\memory[1][0] ),
    .B(_05361_),
    .Y(_07078_)
  );
  OR _15323_ (
    .A(\memory[1][0] ),
    .B(_01491_),
    .Y(_07079_)
  );
  OR _15324_ (
    .A(\data_i[24] ),
    .B(_01492_),
    .Y(_07080_)
  );
  NAND _15325_ (
    .A(_07079_),
    .B(_07080_),
    .Y(_07081_)
  );
  NAND _15326_ (
    .A(_01505_),
    .B(_07081_),
    .Y(_07082_)
  );
  OR _15327_ (
    .A(\data_i[16] ),
    .B(_01505_),
    .Y(_07083_)
  );
  AND _15328_ (
    .A(_07082_),
    .B(_07083_),
    .Y(_07084_)
  );
  NAND _15329_ (
    .A(\data_i[8] ),
    .B(_01449_),
    .Y(_07085_)
  );
  AND _15330_ (
    .A(_01571_),
    .B(_07085_),
    .Y(_07087_)
  );
  NAND _15331_ (
    .A(_01450_),
    .B(_07084_),
    .Y(_07088_)
  );
  NAND _15332_ (
    .A(_07087_),
    .B(_07088_),
    .Y(_07089_)
  );
  OR _15333_ (
    .A(\data_i[0] ),
    .B(_01571_),
    .Y(_07090_)
  );
  AND _15334_ (
    .A(MemWrite_i),
    .B(_07090_),
    .Y(_07091_)
  );
  NAND _15335_ (
    .A(_07089_),
    .B(_07091_),
    .Y(_07092_)
  );
  NAND _15336_ (
    .A(_07078_),
    .B(_07092_),
    .Y(_00088_)
  );
  NAND _15337_ (
    .A(\memory[1][1] ),
    .B(_05361_),
    .Y(_07093_)
  );
  OR _15338_ (
    .A(\memory[1][1] ),
    .B(_01491_),
    .Y(_07094_)
  );
  OR _15339_ (
    .A(\data_i[25] ),
    .B(_01492_),
    .Y(_07095_)
  );
  NAND _15340_ (
    .A(_07094_),
    .B(_07095_),
    .Y(_07097_)
  );
  NAND _15341_ (
    .A(_01505_),
    .B(_07097_),
    .Y(_07098_)
  );
  OR _15342_ (
    .A(\data_i[17] ),
    .B(_01505_),
    .Y(_07099_)
  );
  AND _15343_ (
    .A(_07098_),
    .B(_07099_),
    .Y(_07100_)
  );
  NAND _15344_ (
    .A(\data_i[9] ),
    .B(_01449_),
    .Y(_07101_)
  );
  AND _15345_ (
    .A(_01571_),
    .B(_07101_),
    .Y(_07102_)
  );
  NAND _15346_ (
    .A(_01450_),
    .B(_07100_),
    .Y(_07103_)
  );
  NAND _15347_ (
    .A(_07102_),
    .B(_07103_),
    .Y(_07104_)
  );
  OR _15348_ (
    .A(\data_i[1] ),
    .B(_01571_),
    .Y(_07105_)
  );
  AND _15349_ (
    .A(MemWrite_i),
    .B(_07105_),
    .Y(_07106_)
  );
  NAND _15350_ (
    .A(_07104_),
    .B(_07106_),
    .Y(_07108_)
  );
  NAND _15351_ (
    .A(_07093_),
    .B(_07108_),
    .Y(_00089_)
  );
  NAND _15352_ (
    .A(\memory[1][2] ),
    .B(_05361_),
    .Y(_07109_)
  );
  OR _15353_ (
    .A(\memory[1][2] ),
    .B(_01491_),
    .Y(_07110_)
  );
  OR _15354_ (
    .A(\data_i[26] ),
    .B(_01492_),
    .Y(_07111_)
  );
  NAND _15355_ (
    .A(_07110_),
    .B(_07111_),
    .Y(_07112_)
  );
  NAND _15356_ (
    .A(_01505_),
    .B(_07112_),
    .Y(_07113_)
  );
  OR _15357_ (
    .A(\data_i[18] ),
    .B(_01505_),
    .Y(_07114_)
  );
  AND _15358_ (
    .A(_07113_),
    .B(_07114_),
    .Y(_07115_)
  );
  NAND _15359_ (
    .A(\data_i[10] ),
    .B(_01449_),
    .Y(_07116_)
  );
  AND _15360_ (
    .A(_01571_),
    .B(_07116_),
    .Y(_07118_)
  );
  NAND _15361_ (
    .A(_01450_),
    .B(_07115_),
    .Y(_07119_)
  );
  NAND _15362_ (
    .A(_07118_),
    .B(_07119_),
    .Y(_07120_)
  );
  OR _15363_ (
    .A(\data_i[2] ),
    .B(_01571_),
    .Y(_07121_)
  );
  AND _15364_ (
    .A(MemWrite_i),
    .B(_07121_),
    .Y(_07122_)
  );
  NAND _15365_ (
    .A(_07120_),
    .B(_07122_),
    .Y(_07123_)
  );
  NAND _15366_ (
    .A(_07109_),
    .B(_07123_),
    .Y(_00090_)
  );
  NAND _15367_ (
    .A(\memory[1][3] ),
    .B(_05361_),
    .Y(_07124_)
  );
  OR _15368_ (
    .A(\memory[1][3] ),
    .B(_01491_),
    .Y(_07125_)
  );
  OR _15369_ (
    .A(\data_i[27] ),
    .B(_01492_),
    .Y(_07126_)
  );
  NAND _15370_ (
    .A(_07125_),
    .B(_07126_),
    .Y(_07128_)
  );
  NAND _15371_ (
    .A(_01505_),
    .B(_07128_),
    .Y(_07129_)
  );
  OR _15372_ (
    .A(\data_i[19] ),
    .B(_01505_),
    .Y(_07130_)
  );
  AND _15373_ (
    .A(_07129_),
    .B(_07130_),
    .Y(_07131_)
  );
  NAND _15374_ (
    .A(\data_i[11] ),
    .B(_01449_),
    .Y(_07132_)
  );
  AND _15375_ (
    .A(_01571_),
    .B(_07132_),
    .Y(_07133_)
  );
  NAND _15376_ (
    .A(_01450_),
    .B(_07131_),
    .Y(_07134_)
  );
  NAND _15377_ (
    .A(_07133_),
    .B(_07134_),
    .Y(_07135_)
  );
  OR _15378_ (
    .A(\data_i[3] ),
    .B(_01571_),
    .Y(_07136_)
  );
  AND _15379_ (
    .A(MemWrite_i),
    .B(_07136_),
    .Y(_07137_)
  );
  NAND _15380_ (
    .A(_07135_),
    .B(_07137_),
    .Y(_07139_)
  );
  NAND _15381_ (
    .A(_07124_),
    .B(_07139_),
    .Y(_00091_)
  );
  NAND _15382_ (
    .A(\memory[1][4] ),
    .B(_05361_),
    .Y(_07140_)
  );
  OR _15383_ (
    .A(\memory[1][4] ),
    .B(_01491_),
    .Y(_07141_)
  );
  OR _15384_ (
    .A(\data_i[28] ),
    .B(_01492_),
    .Y(_07142_)
  );
  NAND _15385_ (
    .A(_07141_),
    .B(_07142_),
    .Y(_07143_)
  );
  NAND _15386_ (
    .A(_01505_),
    .B(_07143_),
    .Y(_07144_)
  );
  OR _15387_ (
    .A(\data_i[20] ),
    .B(_01505_),
    .Y(_07145_)
  );
  AND _15388_ (
    .A(_07144_),
    .B(_07145_),
    .Y(_07146_)
  );
  NAND _15389_ (
    .A(\data_i[12] ),
    .B(_01449_),
    .Y(_07147_)
  );
  AND _15390_ (
    .A(_01571_),
    .B(_07147_),
    .Y(_07149_)
  );
  NAND _15391_ (
    .A(_01450_),
    .B(_07146_),
    .Y(_07150_)
  );
  NAND _15392_ (
    .A(_07149_),
    .B(_07150_),
    .Y(_07151_)
  );
  OR _15393_ (
    .A(\data_i[4] ),
    .B(_01571_),
    .Y(_07152_)
  );
  AND _15394_ (
    .A(MemWrite_i),
    .B(_07152_),
    .Y(_07153_)
  );
  NAND _15395_ (
    .A(_07151_),
    .B(_07153_),
    .Y(_07154_)
  );
  NAND _15396_ (
    .A(_07140_),
    .B(_07154_),
    .Y(_00092_)
  );
  NAND _15397_ (
    .A(\memory[1][5] ),
    .B(_05361_),
    .Y(_07155_)
  );
  OR _15398_ (
    .A(\memory[1][5] ),
    .B(_01491_),
    .Y(_07156_)
  );
  OR _15399_ (
    .A(\data_i[29] ),
    .B(_01492_),
    .Y(_07157_)
  );
  NAND _15400_ (
    .A(_07156_),
    .B(_07157_),
    .Y(_07159_)
  );
  NAND _15401_ (
    .A(_01505_),
    .B(_07159_),
    .Y(_07160_)
  );
  OR _15402_ (
    .A(\data_i[21] ),
    .B(_01505_),
    .Y(_07161_)
  );
  AND _15403_ (
    .A(_07160_),
    .B(_07161_),
    .Y(_07162_)
  );
  NAND _15404_ (
    .A(\data_i[13] ),
    .B(_01449_),
    .Y(_07163_)
  );
  AND _15405_ (
    .A(_01571_),
    .B(_07163_),
    .Y(_07164_)
  );
  NAND _15406_ (
    .A(_01450_),
    .B(_07162_),
    .Y(_07165_)
  );
  NAND _15407_ (
    .A(_07164_),
    .B(_07165_),
    .Y(_07166_)
  );
  OR _15408_ (
    .A(\data_i[5] ),
    .B(_01571_),
    .Y(_07167_)
  );
  AND _15409_ (
    .A(MemWrite_i),
    .B(_07167_),
    .Y(_07168_)
  );
  NAND _15410_ (
    .A(_07166_),
    .B(_07168_),
    .Y(_07170_)
  );
  NAND _15411_ (
    .A(_07155_),
    .B(_07170_),
    .Y(_00093_)
  );
  NAND _15412_ (
    .A(\memory[1][6] ),
    .B(_05361_),
    .Y(_07171_)
  );
  OR _15413_ (
    .A(\memory[1][6] ),
    .B(_01491_),
    .Y(_07172_)
  );
  OR _15414_ (
    .A(\data_i[30] ),
    .B(_01492_),
    .Y(_07173_)
  );
  NAND _15415_ (
    .A(_07172_),
    .B(_07173_),
    .Y(_07174_)
  );
  NAND _15416_ (
    .A(_01505_),
    .B(_07174_),
    .Y(_07175_)
  );
  OR _15417_ (
    .A(\data_i[22] ),
    .B(_01505_),
    .Y(_07176_)
  );
  AND _15418_ (
    .A(_07175_),
    .B(_07176_),
    .Y(_07177_)
  );
  NAND _15419_ (
    .A(\data_i[14] ),
    .B(_01449_),
    .Y(_07178_)
  );
  AND _15420_ (
    .A(_01571_),
    .B(_07178_),
    .Y(_07180_)
  );
  NAND _15421_ (
    .A(_01450_),
    .B(_07177_),
    .Y(_07181_)
  );
  NAND _15422_ (
    .A(_07180_),
    .B(_07181_),
    .Y(_07182_)
  );
  OR _15423_ (
    .A(\data_i[6] ),
    .B(_01571_),
    .Y(_07183_)
  );
  AND _15424_ (
    .A(MemWrite_i),
    .B(_07183_),
    .Y(_07184_)
  );
  NAND _15425_ (
    .A(_07182_),
    .B(_07184_),
    .Y(_07185_)
  );
  NAND _15426_ (
    .A(_07171_),
    .B(_07185_),
    .Y(_00094_)
  );
  NAND _15427_ (
    .A(\memory[1][7] ),
    .B(_05361_),
    .Y(_07186_)
  );
  OR _15428_ (
    .A(\memory[1][7] ),
    .B(_01491_),
    .Y(_07187_)
  );
  OR _15429_ (
    .A(\data_i[31] ),
    .B(_01492_),
    .Y(_07188_)
  );
  NAND _15430_ (
    .A(_07187_),
    .B(_07188_),
    .Y(_07190_)
  );
  NAND _15431_ (
    .A(_01505_),
    .B(_07190_),
    .Y(_07191_)
  );
  OR _15432_ (
    .A(\data_i[23] ),
    .B(_01505_),
    .Y(_07192_)
  );
  AND _15433_ (
    .A(_07191_),
    .B(_07192_),
    .Y(_07193_)
  );
  NAND _15434_ (
    .A(\data_i[15] ),
    .B(_01449_),
    .Y(_07194_)
  );
  AND _15435_ (
    .A(_01571_),
    .B(_07194_),
    .Y(_07195_)
  );
  NAND _15436_ (
    .A(_01450_),
    .B(_07193_),
    .Y(_07196_)
  );
  NAND _15437_ (
    .A(_07195_),
    .B(_07196_),
    .Y(_07197_)
  );
  OR _15438_ (
    .A(\data_i[7] ),
    .B(_01571_),
    .Y(_07198_)
  );
  AND _15439_ (
    .A(MemWrite_i),
    .B(_07198_),
    .Y(_07199_)
  );
  NAND _15440_ (
    .A(_07197_),
    .B(_07199_),
    .Y(_07201_)
  );
  NAND _15441_ (
    .A(_07186_),
    .B(_07201_),
    .Y(_00095_)
  );
  NAND _15442_ (
    .A(\memory[0][0] ),
    .B(_05361_),
    .Y(_07202_)
  );
  OR _15443_ (
    .A(\memory[0][0] ),
    .B(_01510_),
    .Y(_07203_)
  );
  OR _15444_ (
    .A(\data_i[24] ),
    .B(_01511_),
    .Y(_07204_)
  );
  NAND _15445_ (
    .A(_07203_),
    .B(_07204_),
    .Y(_07205_)
  );
  NAND _15446_ (
    .A(_01492_),
    .B(_07205_),
    .Y(_07206_)
  );
  OR _15447_ (
    .A(\data_i[16] ),
    .B(_01492_),
    .Y(_07207_)
  );
  AND _15448_ (
    .A(_07206_),
    .B(_07207_),
    .Y(_07208_)
  );
  NAND _15449_ (
    .A(\data_i[8] ),
    .B(_01504_),
    .Y(_07209_)
  );
  AND _15450_ (
    .A(_01450_),
    .B(_07209_),
    .Y(_07211_)
  );
  NAND _15451_ (
    .A(_01505_),
    .B(_07208_),
    .Y(_07212_)
  );
  NAND _15452_ (
    .A(_07211_),
    .B(_07212_),
    .Y(_07213_)
  );
  OR _15453_ (
    .A(\data_i[0] ),
    .B(_01450_),
    .Y(_07214_)
  );
  AND _15454_ (
    .A(MemWrite_i),
    .B(_07214_),
    .Y(_07215_)
  );
  NAND _15455_ (
    .A(_07213_),
    .B(_07215_),
    .Y(_07216_)
  );
  NAND _15456_ (
    .A(_07202_),
    .B(_07216_),
    .Y(_00000_)
  );
  NAND _15457_ (
    .A(\memory[0][1] ),
    .B(_05361_),
    .Y(_07217_)
  );
  OR _15458_ (
    .A(\memory[0][1] ),
    .B(_01510_),
    .Y(_07218_)
  );
  OR _15459_ (
    .A(\data_i[25] ),
    .B(_01511_),
    .Y(_07219_)
  );
  NAND _15460_ (
    .A(_07218_),
    .B(_07219_),
    .Y(_07221_)
  );
  NAND _15461_ (
    .A(_01492_),
    .B(_07221_),
    .Y(_07222_)
  );
  OR _15462_ (
    .A(\data_i[17] ),
    .B(_01492_),
    .Y(_07223_)
  );
  AND _15463_ (
    .A(_07222_),
    .B(_07223_),
    .Y(_07224_)
  );
  NAND _15464_ (
    .A(\data_i[9] ),
    .B(_01504_),
    .Y(_07225_)
  );
  AND _15465_ (
    .A(_01450_),
    .B(_07225_),
    .Y(_07226_)
  );
  NAND _15466_ (
    .A(_01505_),
    .B(_07224_),
    .Y(_07227_)
  );
  NAND _15467_ (
    .A(_07226_),
    .B(_07227_),
    .Y(_07228_)
  );
  OR _15468_ (
    .A(\data_i[1] ),
    .B(_01450_),
    .Y(_07229_)
  );
  AND _15469_ (
    .A(MemWrite_i),
    .B(_07229_),
    .Y(_07230_)
  );
  NAND _15470_ (
    .A(_07228_),
    .B(_07230_),
    .Y(_07232_)
  );
  NAND _15471_ (
    .A(_07217_),
    .B(_07232_),
    .Y(_00001_)
  );
  NAND _15472_ (
    .A(\memory[0][2] ),
    .B(_05361_),
    .Y(_07233_)
  );
  OR _15473_ (
    .A(\memory[0][2] ),
    .B(_01510_),
    .Y(_07234_)
  );
  OR _15474_ (
    .A(\data_i[26] ),
    .B(_01511_),
    .Y(_07235_)
  );
  NAND _15475_ (
    .A(_07234_),
    .B(_07235_),
    .Y(_07236_)
  );
  NAND _15476_ (
    .A(_01492_),
    .B(_07236_),
    .Y(_07237_)
  );
  OR _15477_ (
    .A(\data_i[18] ),
    .B(_01492_),
    .Y(_07238_)
  );
  AND _15478_ (
    .A(_07237_),
    .B(_07238_),
    .Y(_07239_)
  );
  NAND _15479_ (
    .A(\data_i[10] ),
    .B(_01504_),
    .Y(_07240_)
  );
  AND _15480_ (
    .A(_01450_),
    .B(_07240_),
    .Y(_07242_)
  );
  NAND _15481_ (
    .A(_01505_),
    .B(_07239_),
    .Y(_07243_)
  );
  NAND _15482_ (
    .A(_07242_),
    .B(_07243_),
    .Y(_07244_)
  );
  OR _15483_ (
    .A(\data_i[2] ),
    .B(_01450_),
    .Y(_07245_)
  );
  AND _15484_ (
    .A(MemWrite_i),
    .B(_07245_),
    .Y(_07246_)
  );
  NAND _15485_ (
    .A(_07244_),
    .B(_07246_),
    .Y(_07247_)
  );
  NAND _15486_ (
    .A(_07233_),
    .B(_07247_),
    .Y(_00002_)
  );
  NAND _15487_ (
    .A(\memory[0][3] ),
    .B(_05361_),
    .Y(_07248_)
  );
  OR _15488_ (
    .A(\memory[0][3] ),
    .B(_01510_),
    .Y(_07249_)
  );
  OR _15489_ (
    .A(\data_i[27] ),
    .B(_01511_),
    .Y(_07250_)
  );
  NAND _15490_ (
    .A(_07249_),
    .B(_07250_),
    .Y(_07252_)
  );
  NAND _15491_ (
    .A(_01492_),
    .B(_07252_),
    .Y(_07253_)
  );
  OR _15492_ (
    .A(\data_i[19] ),
    .B(_01492_),
    .Y(_07254_)
  );
  AND _15493_ (
    .A(_07253_),
    .B(_07254_),
    .Y(_07255_)
  );
  NAND _15494_ (
    .A(\data_i[11] ),
    .B(_01504_),
    .Y(_07256_)
  );
  AND _15495_ (
    .A(_01450_),
    .B(_07256_),
    .Y(_07257_)
  );
  NAND _15496_ (
    .A(_01505_),
    .B(_07255_),
    .Y(_07258_)
  );
  NAND _15497_ (
    .A(_07257_),
    .B(_07258_),
    .Y(_07259_)
  );
  OR _15498_ (
    .A(\data_i[3] ),
    .B(_01450_),
    .Y(_07260_)
  );
  AND _15499_ (
    .A(MemWrite_i),
    .B(_07260_),
    .Y(_07261_)
  );
  NAND _15500_ (
    .A(_07259_),
    .B(_07261_),
    .Y(_07263_)
  );
  NAND _15501_ (
    .A(_07248_),
    .B(_07263_),
    .Y(_00003_)
  );
  NAND _15502_ (
    .A(\memory[0][4] ),
    .B(_05361_),
    .Y(_07264_)
  );
  OR _15503_ (
    .A(\memory[0][4] ),
    .B(_01510_),
    .Y(_07265_)
  );
  OR _15504_ (
    .A(\data_i[28] ),
    .B(_01511_),
    .Y(_07266_)
  );
  NAND _15505_ (
    .A(_07265_),
    .B(_07266_),
    .Y(_07267_)
  );
  NAND _15506_ (
    .A(_01492_),
    .B(_07267_),
    .Y(_07268_)
  );
  OR _15507_ (
    .A(\data_i[20] ),
    .B(_01492_),
    .Y(_07269_)
  );
  AND _15508_ (
    .A(_07268_),
    .B(_07269_),
    .Y(_07270_)
  );
  NAND _15509_ (
    .A(\data_i[12] ),
    .B(_01504_),
    .Y(_07271_)
  );
  AND _15510_ (
    .A(_01450_),
    .B(_07271_),
    .Y(_07273_)
  );
  NAND _15511_ (
    .A(_01505_),
    .B(_07270_),
    .Y(_07274_)
  );
  NAND _15512_ (
    .A(_07273_),
    .B(_07274_),
    .Y(_07275_)
  );
  OR _15513_ (
    .A(\data_i[4] ),
    .B(_01450_),
    .Y(_07276_)
  );
  AND _15514_ (
    .A(MemWrite_i),
    .B(_07276_),
    .Y(_07277_)
  );
  NAND _15515_ (
    .A(_07275_),
    .B(_07277_),
    .Y(_07278_)
  );
  NAND _15516_ (
    .A(_07264_),
    .B(_07278_),
    .Y(_00004_)
  );
  NAND _15517_ (
    .A(\memory[0][5] ),
    .B(_05361_),
    .Y(_07279_)
  );
  OR _15518_ (
    .A(\memory[0][5] ),
    .B(_01510_),
    .Y(_07280_)
  );
  OR _15519_ (
    .A(\data_i[29] ),
    .B(_01511_),
    .Y(_07281_)
  );
  NAND _15520_ (
    .A(_07280_),
    .B(_07281_),
    .Y(_07283_)
  );
  NAND _15521_ (
    .A(_01492_),
    .B(_07283_),
    .Y(_07284_)
  );
  OR _15522_ (
    .A(\data_i[21] ),
    .B(_01492_),
    .Y(_07285_)
  );
  AND _15523_ (
    .A(_07284_),
    .B(_07285_),
    .Y(_07286_)
  );
  NAND _15524_ (
    .A(\data_i[13] ),
    .B(_01504_),
    .Y(_07287_)
  );
  AND _15525_ (
    .A(_01450_),
    .B(_07287_),
    .Y(_07288_)
  );
  NAND _15526_ (
    .A(_01505_),
    .B(_07286_),
    .Y(_07289_)
  );
  NAND _15527_ (
    .A(_07288_),
    .B(_07289_),
    .Y(_07290_)
  );
  OR _15528_ (
    .A(\data_i[5] ),
    .B(_01450_),
    .Y(_07291_)
  );
  AND _15529_ (
    .A(MemWrite_i),
    .B(_07291_),
    .Y(_07292_)
  );
  NAND _15530_ (
    .A(_07290_),
    .B(_07292_),
    .Y(_07294_)
  );
  NAND _15531_ (
    .A(_07279_),
    .B(_07294_),
    .Y(_00005_)
  );
  NAND _15532_ (
    .A(\memory[0][6] ),
    .B(_05361_),
    .Y(_07295_)
  );
  OR _15533_ (
    .A(\memory[0][6] ),
    .B(_01510_),
    .Y(_07296_)
  );
  OR _15534_ (
    .A(\data_i[30] ),
    .B(_01511_),
    .Y(_07297_)
  );
  NAND _15535_ (
    .A(_07296_),
    .B(_07297_),
    .Y(_07298_)
  );
  NAND _15536_ (
    .A(_01492_),
    .B(_07298_),
    .Y(_07299_)
  );
  OR _15537_ (
    .A(\data_i[22] ),
    .B(_01492_),
    .Y(_07300_)
  );
  AND _15538_ (
    .A(_07299_),
    .B(_07300_),
    .Y(_07301_)
  );
  NAND _15539_ (
    .A(\data_i[14] ),
    .B(_01504_),
    .Y(_07302_)
  );
  AND _15540_ (
    .A(_01450_),
    .B(_07302_),
    .Y(_07304_)
  );
  NAND _15541_ (
    .A(_01505_),
    .B(_07301_),
    .Y(_07305_)
  );
  NAND _15542_ (
    .A(_07304_),
    .B(_07305_),
    .Y(_07306_)
  );
  OR _15543_ (
    .A(\data_i[6] ),
    .B(_01450_),
    .Y(_07307_)
  );
  AND _15544_ (
    .A(MemWrite_i),
    .B(_07307_),
    .Y(_07308_)
  );
  NAND _15545_ (
    .A(_07306_),
    .B(_07308_),
    .Y(_07309_)
  );
  NAND _15546_ (
    .A(_07295_),
    .B(_07309_),
    .Y(_00006_)
  );
  NAND _15547_ (
    .A(\memory[0][7] ),
    .B(_05361_),
    .Y(_07310_)
  );
  OR _15548_ (
    .A(\memory[0][7] ),
    .B(_01510_),
    .Y(_07311_)
  );
  OR _15549_ (
    .A(\data_i[31] ),
    .B(_01511_),
    .Y(_07312_)
  );
  NAND _15550_ (
    .A(_07311_),
    .B(_07312_),
    .Y(_07314_)
  );
  NAND _15551_ (
    .A(_01492_),
    .B(_07314_),
    .Y(_07315_)
  );
  OR _15552_ (
    .A(\data_i[23] ),
    .B(_01492_),
    .Y(_07316_)
  );
  AND _15553_ (
    .A(_07315_),
    .B(_07316_),
    .Y(_07317_)
  );
  NAND _15554_ (
    .A(\data_i[15] ),
    .B(_01504_),
    .Y(_07318_)
  );
  AND _15555_ (
    .A(_01450_),
    .B(_07318_),
    .Y(_07319_)
  );
  NAND _15556_ (
    .A(_01505_),
    .B(_07317_),
    .Y(_07320_)
  );
  NAND _15557_ (
    .A(_07319_),
    .B(_07320_),
    .Y(_07321_)
  );
  OR _15558_ (
    .A(\data_i[7] ),
    .B(_01450_),
    .Y(_07322_)
  );
  AND _15559_ (
    .A(MemWrite_i),
    .B(_07322_),
    .Y(_07323_)
  );
  NAND _15560_ (
    .A(_07321_),
    .B(_07323_),
    .Y(_07325_)
  );
  NAND _15561_ (
    .A(_07310_),
    .B(_07325_),
    .Y(_00007_)
  );
  NAND _15562_ (
    .A(\memory[30][0] ),
    .B(_05847_),
    .Y(_07326_)
  );
  NAND _15563_ (
    .A(\memory[14][0] ),
    .B(_05785_),
    .Y(_07327_)
  );
  NAND _15564_ (
    .A(\memory[7][0] ),
    .B(_05733_),
    .Y(_07328_)
  );
  NAND _15565_ (
    .A(\memory[19][0] ),
    .B(_05558_),
    .Y(_07329_)
  );
  NAND _15566_ (
    .A(\memory[15][0] ),
    .B(_06002_),
    .Y(_07330_)
  );
  NAND _15567_ (
    .A(\memory[13][0] ),
    .B(_05661_),
    .Y(_07331_)
  );
  NAND _15568_ (
    .A(\memory[23][0] ),
    .B(_05806_),
    .Y(_07332_)
  );
  NAND _15569_ (
    .A(\memory[24][0] ),
    .B(_06023_),
    .Y(_07333_)
  );
  NAND _15570_ (
    .A(\memory[3][0] ),
    .B(_06043_),
    .Y(_07335_)
  );
  NAND _15571_ (
    .A(\memory[8][0] ),
    .B(_05475_),
    .Y(_07336_)
  );
  NAND _15572_ (
    .A(\memory[16][0] ),
    .B(_06064_),
    .Y(_07337_)
  );
  NAND _15573_ (
    .A(\memory[12][0] ),
    .B(_06312_),
    .Y(_07338_)
  );
  NAND _15574_ (
    .A(\memory[10][0] ),
    .B(_06353_),
    .Y(_07339_)
  );
  NAND _15575_ (
    .A(\memory[27][0] ),
    .B(_06333_),
    .Y(_07340_)
  );
  NAND _15576_ (
    .A(\memory[29][0] ),
    .B(_05981_),
    .Y(_07341_)
  );
  NAND _15577_ (
    .A(\memory[31][0] ),
    .B(_05826_),
    .Y(_07342_)
  );
  NAND _15578_ (
    .A(\memory[0][0] ),
    .B(_05692_),
    .Y(_07343_)
  );
  AND _15579_ (
    .A(_07342_),
    .B(_07343_),
    .Y(_07344_)
  );
  NAND _15580_ (
    .A(\memory[4][0] ),
    .B(_05599_),
    .Y(_07346_)
  );
  NAND _15581_ (
    .A(\memory[20][0] ),
    .B(_05754_),
    .Y(_07347_)
  );
  NAND _15582_ (
    .A(\memory[28][0] ),
    .B(_06291_),
    .Y(_07348_)
  );
  NAND _15583_ (
    .A(\memory[1][0] ),
    .B(_06188_),
    .Y(_07349_)
  );
  NAND _15584_ (
    .A(\memory[6][0] ),
    .B(_06147_),
    .Y(_07350_)
  );
  NAND _15585_ (
    .A(\memory[22][0] ),
    .B(_06167_),
    .Y(_07351_)
  );
  NAND _15586_ (
    .A(\memory[2][0] ),
    .B(_06116_),
    .Y(_07352_)
  );
  NAND _15587_ (
    .A(\memory[18][0] ),
    .B(_06209_),
    .Y(_07353_)
  );
  NAND _15588_ (
    .A(\memory[21][0] ),
    .B(_05930_),
    .Y(_07354_)
  );
  NAND _15589_ (
    .A(\memory[25][0] ),
    .B(_06395_),
    .Y(_07355_)
  );
  NAND _15590_ (
    .A(\memory[9][0] ),
    .B(_06374_),
    .Y(_07357_)
  );
  NAND _15591_ (
    .A(\memory[5][0] ),
    .B(_05961_),
    .Y(_07358_)
  );
  NAND _15592_ (
    .A(\memory[11][0] ),
    .B(_05899_),
    .Y(_07359_)
  );
  NAND _15593_ (
    .A(\memory[17][0] ),
    .B(_06085_),
    .Y(_07360_)
  );
  NAND _15594_ (
    .A(\memory[26][0] ),
    .B(_06250_),
    .Y(_07361_)
  );
  AND _15595_ (
    .A(_07355_),
    .B(_07361_),
    .Y(_07362_)
  );
  AND _15596_ (
    .A(_07341_),
    .B(_07360_),
    .Y(_07363_)
  );
  AND _15597_ (
    .A(_07350_),
    .B(_07358_),
    .Y(_07364_)
  );
  AND _15598_ (
    .A(_07346_),
    .B(_07364_),
    .Y(_07365_)
  );
  AND _15599_ (
    .A(_07331_),
    .B(_07359_),
    .Y(_07366_)
  );
  AND _15600_ (
    .A(_07340_),
    .B(_07354_),
    .Y(_07368_)
  );
  AND _15601_ (
    .A(_07366_),
    .B(_07368_),
    .Y(_07369_)
  );
  AND _15602_ (
    .A(_07349_),
    .B(_07369_),
    .Y(_07370_)
  );
  AND _15603_ (
    .A(_07327_),
    .B(_07338_),
    .Y(_07371_)
  );
  AND _15604_ (
    .A(_07363_),
    .B(_07371_),
    .Y(_07372_)
  );
  AND _15605_ (
    .A(_07328_),
    .B(_07336_),
    .Y(_07373_)
  );
  AND _15606_ (
    .A(_07352_),
    .B(_07373_),
    .Y(_07374_)
  );
  AND _15607_ (
    .A(_07339_),
    .B(_07374_),
    .Y(_07375_)
  );
  AND _15608_ (
    .A(_07372_),
    .B(_07375_),
    .Y(_07376_)
  );
  AND _15609_ (
    .A(_07370_),
    .B(_07376_),
    .Y(_07377_)
  );
  AND _15610_ (
    .A(_07333_),
    .B(_07347_),
    .Y(_07378_)
  );
  AND _15611_ (
    .A(_07332_),
    .B(_07351_),
    .Y(_07379_)
  );
  AND _15612_ (
    .A(_07326_),
    .B(_07379_),
    .Y(_07380_)
  );
  AND _15613_ (
    .A(_07378_),
    .B(_07380_),
    .Y(_07381_)
  );
  AND _15614_ (
    .A(_07344_),
    .B(_07362_),
    .Y(_07382_)
  );
  AND _15615_ (
    .A(_07381_),
    .B(_07382_),
    .Y(_07383_)
  );
  AND _15616_ (
    .A(_07329_),
    .B(_07348_),
    .Y(_07384_)
  );
  AND _15617_ (
    .A(_07353_),
    .B(_07384_),
    .Y(_07385_)
  );
  AND _15618_ (
    .A(_07330_),
    .B(_07337_),
    .Y(_07386_)
  );
  AND _15619_ (
    .A(_07335_),
    .B(_07357_),
    .Y(_07387_)
  );
  AND _15620_ (
    .A(_07386_),
    .B(_07387_),
    .Y(_07389_)
  );
  AND _15621_ (
    .A(_07385_),
    .B(_07389_),
    .Y(_07390_)
  );
  AND _15622_ (
    .A(_07383_),
    .B(_07390_),
    .Y(_07391_)
  );
  AND _15623_ (
    .A(_07377_),
    .B(_07391_),
    .Y(_07392_)
  );
  NAND _15624_ (
    .A(_07365_),
    .B(_07392_),
    .Y(\data_mem_o[24] )
  );
  NAND _15625_ (
    .A(\memory[20][1] ),
    .B(_05754_),
    .Y(_07393_)
  );
  NAND _15626_ (
    .A(\memory[16][1] ),
    .B(_06064_),
    .Y(_07394_)
  );
  NAND _15627_ (
    .A(\memory[3][1] ),
    .B(_06043_),
    .Y(_07395_)
  );
  NAND _15628_ (
    .A(\memory[31][1] ),
    .B(_05826_),
    .Y(_07396_)
  );
  NAND _15629_ (
    .A(\memory[0][1] ),
    .B(_05692_),
    .Y(_07397_)
  );
  AND _15630_ (
    .A(_07396_),
    .B(_07397_),
    .Y(_07399_)
  );
  NAND _15631_ (
    .A(\memory[4][1] ),
    .B(_05599_),
    .Y(_07400_)
  );
  NAND _15632_ (
    .A(\memory[30][1] ),
    .B(_05847_),
    .Y(_07401_)
  );
  NAND _15633_ (
    .A(\memory[7][1] ),
    .B(_05733_),
    .Y(_07402_)
  );
  NAND _15634_ (
    .A(\memory[15][1] ),
    .B(_06002_),
    .Y(_07403_)
  );
  NAND _15635_ (
    .A(\memory[14][1] ),
    .B(_05785_),
    .Y(_07404_)
  );
  NAND _15636_ (
    .A(\memory[24][1] ),
    .B(_06023_),
    .Y(_07405_)
  );
  NAND _15637_ (
    .A(\memory[12][1] ),
    .B(_06312_),
    .Y(_07406_)
  );
  NAND _15638_ (
    .A(\memory[10][1] ),
    .B(_06353_),
    .Y(_07407_)
  );
  NAND _15639_ (
    .A(\memory[27][1] ),
    .B(_06333_),
    .Y(_07408_)
  );
  NAND _15640_ (
    .A(\memory[29][1] ),
    .B(_05981_),
    .Y(_07410_)
  );
  NAND _15641_ (
    .A(\memory[13][1] ),
    .B(_05661_),
    .Y(_07411_)
  );
  NAND _15642_ (
    .A(\memory[8][1] ),
    .B(_05475_),
    .Y(_07412_)
  );
  NAND _15643_ (
    .A(\memory[23][1] ),
    .B(_05806_),
    .Y(_07413_)
  );
  NAND _15644_ (
    .A(\memory[19][1] ),
    .B(_05558_),
    .Y(_07414_)
  );
  NAND _15645_ (
    .A(\memory[28][1] ),
    .B(_06291_),
    .Y(_07415_)
  );
  NAND _15646_ (
    .A(\memory[1][1] ),
    .B(_06188_),
    .Y(_07416_)
  );
  NAND _15647_ (
    .A(\memory[18][1] ),
    .B(_06209_),
    .Y(_07417_)
  );
  NAND _15648_ (
    .A(\memory[2][1] ),
    .B(_06116_),
    .Y(_07418_)
  );
  NAND _15649_ (
    .A(\memory[6][1] ),
    .B(_06147_),
    .Y(_07419_)
  );
  NAND _15650_ (
    .A(\memory[22][1] ),
    .B(_06167_),
    .Y(_07421_)
  );
  NAND _15651_ (
    .A(\memory[9][1] ),
    .B(_06374_),
    .Y(_07422_)
  );
  NAND _15652_ (
    .A(\memory[11][1] ),
    .B(_05899_),
    .Y(_07423_)
  );
  NAND _15653_ (
    .A(\memory[25][1] ),
    .B(_06395_),
    .Y(_07424_)
  );
  NAND _15654_ (
    .A(\memory[21][1] ),
    .B(_05930_),
    .Y(_07425_)
  );
  NAND _15655_ (
    .A(\memory[17][1] ),
    .B(_06085_),
    .Y(_07426_)
  );
  NAND _15656_ (
    .A(\memory[5][1] ),
    .B(_05961_),
    .Y(_07427_)
  );
  NAND _15657_ (
    .A(\memory[26][1] ),
    .B(_06250_),
    .Y(_07428_)
  );
  AND _15658_ (
    .A(_07424_),
    .B(_07428_),
    .Y(_07429_)
  );
  AND _15659_ (
    .A(_07410_),
    .B(_07426_),
    .Y(_07430_)
  );
  AND _15660_ (
    .A(_07419_),
    .B(_07427_),
    .Y(_07432_)
  );
  AND _15661_ (
    .A(_07400_),
    .B(_07432_),
    .Y(_07433_)
  );
  AND _15662_ (
    .A(_07411_),
    .B(_07423_),
    .Y(_07434_)
  );
  AND _15663_ (
    .A(_07408_),
    .B(_07425_),
    .Y(_07435_)
  );
  AND _15664_ (
    .A(_07434_),
    .B(_07435_),
    .Y(_07436_)
  );
  AND _15665_ (
    .A(_07416_),
    .B(_07436_),
    .Y(_07437_)
  );
  AND _15666_ (
    .A(_07404_),
    .B(_07406_),
    .Y(_07438_)
  );
  AND _15667_ (
    .A(_07430_),
    .B(_07438_),
    .Y(_07439_)
  );
  AND _15668_ (
    .A(_07402_),
    .B(_07412_),
    .Y(_07440_)
  );
  AND _15669_ (
    .A(_07418_),
    .B(_07440_),
    .Y(_07441_)
  );
  AND _15670_ (
    .A(_07407_),
    .B(_07441_),
    .Y(_07443_)
  );
  AND _15671_ (
    .A(_07439_),
    .B(_07443_),
    .Y(_07444_)
  );
  AND _15672_ (
    .A(_07437_),
    .B(_07444_),
    .Y(_07445_)
  );
  AND _15673_ (
    .A(_07393_),
    .B(_07405_),
    .Y(_07446_)
  );
  AND _15674_ (
    .A(_07413_),
    .B(_07421_),
    .Y(_07447_)
  );
  AND _15675_ (
    .A(_07401_),
    .B(_07447_),
    .Y(_07448_)
  );
  AND _15676_ (
    .A(_07446_),
    .B(_07448_),
    .Y(_07449_)
  );
  AND _15677_ (
    .A(_07399_),
    .B(_07429_),
    .Y(_07450_)
  );
  AND _15678_ (
    .A(_07449_),
    .B(_07450_),
    .Y(_07451_)
  );
  AND _15679_ (
    .A(_07414_),
    .B(_07415_),
    .Y(_07452_)
  );
  AND _15680_ (
    .A(_07417_),
    .B(_07452_),
    .Y(_07454_)
  );
  AND _15681_ (
    .A(_07394_),
    .B(_07403_),
    .Y(_07455_)
  );
  AND _15682_ (
    .A(_07395_),
    .B(_07422_),
    .Y(_07456_)
  );
  AND _15683_ (
    .A(_07455_),
    .B(_07456_),
    .Y(_07457_)
  );
  AND _15684_ (
    .A(_07454_),
    .B(_07457_),
    .Y(_07458_)
  );
  AND _15685_ (
    .A(_07451_),
    .B(_07458_),
    .Y(_07459_)
  );
  AND _15686_ (
    .A(_07445_),
    .B(_07459_),
    .Y(_07460_)
  );
  NAND _15687_ (
    .A(_07433_),
    .B(_07460_),
    .Y(\data_mem_o[25] )
  );
  NAND _15688_ (
    .A(\memory[3][2] ),
    .B(_06043_),
    .Y(_07461_)
  );
  NAND _15689_ (
    .A(\memory[16][2] ),
    .B(_06064_),
    .Y(_07462_)
  );
  NAND _15690_ (
    .A(\memory[23][2] ),
    .B(_05806_),
    .Y(_07464_)
  );
  NAND _15691_ (
    .A(\memory[24][2] ),
    .B(_06023_),
    .Y(_07465_)
  );
  NAND _15692_ (
    .A(\memory[31][2] ),
    .B(_05826_),
    .Y(_07466_)
  );
  NAND _15693_ (
    .A(\memory[20][2] ),
    .B(_05754_),
    .Y(_07467_)
  );
  NAND _15694_ (
    .A(\memory[4][2] ),
    .B(_05599_),
    .Y(_07468_)
  );
  NAND _15695_ (
    .A(\memory[14][2] ),
    .B(_05785_),
    .Y(_07469_)
  );
  NAND _15696_ (
    .A(\memory[30][2] ),
    .B(_05847_),
    .Y(_07470_)
  );
  NAND _15697_ (
    .A(\memory[15][2] ),
    .B(_06002_),
    .Y(_07471_)
  );
  NAND _15698_ (
    .A(\memory[0][2] ),
    .B(_05692_),
    .Y(_07472_)
  );
  NAND _15699_ (
    .A(\memory[9][2] ),
    .B(_06374_),
    .Y(_07473_)
  );
  NAND _15700_ (
    .A(\memory[29][2] ),
    .B(_05981_),
    .Y(_07475_)
  );
  NAND _15701_ (
    .A(\memory[17][2] ),
    .B(_06085_),
    .Y(_07476_)
  );
  NAND _15702_ (
    .A(\memory[21][2] ),
    .B(_05930_),
    .Y(_07477_)
  );
  NAND _15703_ (
    .A(\memory[13][2] ),
    .B(_05661_),
    .Y(_07478_)
  );
  NAND _15704_ (
    .A(\memory[19][2] ),
    .B(_05558_),
    .Y(_07479_)
  );
  NAND _15705_ (
    .A(\memory[7][2] ),
    .B(_05733_),
    .Y(_07480_)
  );
  NAND _15706_ (
    .A(\memory[8][2] ),
    .B(_05475_),
    .Y(_07481_)
  );
  NAND _15707_ (
    .A(\memory[25][2] ),
    .B(_06395_),
    .Y(_07482_)
  );
  NAND _15708_ (
    .A(\memory[1][2] ),
    .B(_06188_),
    .Y(_07483_)
  );
  NAND _15709_ (
    .A(\memory[22][2] ),
    .B(_06167_),
    .Y(_07484_)
  );
  NAND _15710_ (
    .A(\memory[6][2] ),
    .B(_06147_),
    .Y(_07486_)
  );
  NAND _15711_ (
    .A(\memory[2][2] ),
    .B(_06116_),
    .Y(_07487_)
  );
  NAND _15712_ (
    .A(\memory[18][2] ),
    .B(_06209_),
    .Y(_07488_)
  );
  NAND _15713_ (
    .A(\memory[12][2] ),
    .B(_06312_),
    .Y(_07489_)
  );
  NAND _15714_ (
    .A(\memory[10][2] ),
    .B(_06353_),
    .Y(_07490_)
  );
  NAND _15715_ (
    .A(\memory[28][2] ),
    .B(_06291_),
    .Y(_07491_)
  );
  NAND _15716_ (
    .A(\memory[26][2] ),
    .B(_06250_),
    .Y(_07492_)
  );
  NAND _15717_ (
    .A(\memory[27][2] ),
    .B(_06333_),
    .Y(_07493_)
  );
  AND _15718_ (
    .A(_07492_),
    .B(_07493_),
    .Y(_07494_)
  );
  NAND _15719_ (
    .A(\memory[5][2] ),
    .B(_05961_),
    .Y(_07495_)
  );
  NAND _15720_ (
    .A(\memory[11][2] ),
    .B(_05899_),
    .Y(_07497_)
  );
  AND _15721_ (
    .A(_07468_),
    .B(_07495_),
    .Y(_07498_)
  );
  AND _15722_ (
    .A(_07478_),
    .B(_07483_),
    .Y(_07499_)
  );
  AND _15723_ (
    .A(_07461_),
    .B(_07489_),
    .Y(_07500_)
  );
  AND _15724_ (
    .A(_07498_),
    .B(_07500_),
    .Y(_07501_)
  );
  AND _15725_ (
    .A(_07499_),
    .B(_07501_),
    .Y(_07502_)
  );
  AND _15726_ (
    .A(_07467_),
    .B(_07502_),
    .Y(_07503_)
  );
  AND _15727_ (
    .A(_07469_),
    .B(_07487_),
    .Y(_07504_)
  );
  AND _15728_ (
    .A(_07484_),
    .B(_07488_),
    .Y(_07505_)
  );
  AND _15729_ (
    .A(_07462_),
    .B(_07505_),
    .Y(_07506_)
  );
  AND _15730_ (
    .A(_07464_),
    .B(_07465_),
    .Y(_07508_)
  );
  AND _15731_ (
    .A(_07471_),
    .B(_07508_),
    .Y(_07509_)
  );
  AND _15732_ (
    .A(_07506_),
    .B(_07509_),
    .Y(_07510_)
  );
  AND _15733_ (
    .A(_07476_),
    .B(_07479_),
    .Y(_07511_)
  );
  AND _15734_ (
    .A(_07477_),
    .B(_07482_),
    .Y(_07512_)
  );
  AND _15735_ (
    .A(_07511_),
    .B(_07512_),
    .Y(_07513_)
  );
  AND _15736_ (
    .A(_07510_),
    .B(_07513_),
    .Y(_07514_)
  );
  AND _15737_ (
    .A(_07504_),
    .B(_07514_),
    .Y(_07515_)
  );
  AND _15738_ (
    .A(_07503_),
    .B(_07515_),
    .Y(_07516_)
  );
  AND _15739_ (
    .A(_07466_),
    .B(_07470_),
    .Y(_07517_)
  );
  AND _15740_ (
    .A(_07480_),
    .B(_07490_),
    .Y(_07519_)
  );
  AND _15741_ (
    .A(_07517_),
    .B(_07519_),
    .Y(_07520_)
  );
  AND _15742_ (
    .A(_07486_),
    .B(_07497_),
    .Y(_07521_)
  );
  AND _15743_ (
    .A(_07473_),
    .B(_07521_),
    .Y(_07522_)
  );
  AND _15744_ (
    .A(_07472_),
    .B(_07475_),
    .Y(_07523_)
  );
  AND _15745_ (
    .A(_07481_),
    .B(_07491_),
    .Y(_07524_)
  );
  AND _15746_ (
    .A(_07523_),
    .B(_07524_),
    .Y(_07525_)
  );
  AND _15747_ (
    .A(_07522_),
    .B(_07525_),
    .Y(_07526_)
  );
  AND _15748_ (
    .A(_07494_),
    .B(_07526_),
    .Y(_07527_)
  );
  AND _15749_ (
    .A(_07520_),
    .B(_07527_),
    .Y(_07528_)
  );
  NAND _15750_ (
    .A(_07516_),
    .B(_07528_),
    .Y(\data_mem_o[26] )
  );
  NAND _15751_ (
    .A(\memory[4][3] ),
    .B(_05599_),
    .Y(_07530_)
  );
  NAND _15752_ (
    .A(\memory[30][3] ),
    .B(_05847_),
    .Y(_07531_)
  );
  NAND _15753_ (
    .A(\memory[8][3] ),
    .B(_05475_),
    .Y(_07532_)
  );
  NAND _15754_ (
    .A(\memory[31][3] ),
    .B(_05826_),
    .Y(_07533_)
  );
  NAND _15755_ (
    .A(\memory[0][3] ),
    .B(_05692_),
    .Y(_07534_)
  );
  NAND _15756_ (
    .A(\memory[20][3] ),
    .B(_05754_),
    .Y(_07535_)
  );
  NAND _15757_ (
    .A(\memory[7][3] ),
    .B(_05733_),
    .Y(_07536_)
  );
  NAND _15758_ (
    .A(\memory[23][3] ),
    .B(_05806_),
    .Y(_07537_)
  );
  NAND _15759_ (
    .A(\memory[16][3] ),
    .B(_06064_),
    .Y(_07538_)
  );
  NAND _15760_ (
    .A(\memory[3][3] ),
    .B(_06043_),
    .Y(_07540_)
  );
  NAND _15761_ (
    .A(\memory[19][3] ),
    .B(_05558_),
    .Y(_07541_)
  );
  NAND _15762_ (
    .A(\memory[17][3] ),
    .B(_06085_),
    .Y(_07542_)
  );
  NAND _15763_ (
    .A(\memory[29][3] ),
    .B(_05981_),
    .Y(_07543_)
  );
  NAND _15764_ (
    .A(\memory[9][3] ),
    .B(_06374_),
    .Y(_07544_)
  );
  NAND _15765_ (
    .A(\memory[26][3] ),
    .B(_06250_),
    .Y(_07545_)
  );
  NAND _15766_ (
    .A(\memory[14][3] ),
    .B(_05785_),
    .Y(_07546_)
  );
  NAND _15767_ (
    .A(\memory[24][3] ),
    .B(_06023_),
    .Y(_07547_)
  );
  NAND _15768_ (
    .A(\memory[13][3] ),
    .B(_05661_),
    .Y(_07548_)
  );
  NAND _15769_ (
    .A(\memory[15][3] ),
    .B(_06002_),
    .Y(_07549_)
  );
  NAND _15770_ (
    .A(\memory[5][3] ),
    .B(_05961_),
    .Y(_07551_)
  );
  NAND _15771_ (
    .A(\memory[18][3] ),
    .B(_06209_),
    .Y(_07552_)
  );
  NAND _15772_ (
    .A(\memory[6][3] ),
    .B(_06147_),
    .Y(_07553_)
  );
  NAND _15773_ (
    .A(\memory[22][3] ),
    .B(_06167_),
    .Y(_07554_)
  );
  NAND _15774_ (
    .A(\memory[2][3] ),
    .B(_06116_),
    .Y(_07555_)
  );
  NAND _15775_ (
    .A(\memory[1][3] ),
    .B(_06188_),
    .Y(_07556_)
  );
  NAND _15776_ (
    .A(\memory[11][3] ),
    .B(_05899_),
    .Y(_07557_)
  );
  NAND _15777_ (
    .A(\memory[25][3] ),
    .B(_06395_),
    .Y(_07558_)
  );
  NAND _15778_ (
    .A(\memory[28][3] ),
    .B(_06291_),
    .Y(_07559_)
  );
  NAND _15779_ (
    .A(\memory[21][3] ),
    .B(_05930_),
    .Y(_07560_)
  );
  NAND _15780_ (
    .A(\memory[10][3] ),
    .B(_06353_),
    .Y(_07562_)
  );
  NAND _15781_ (
    .A(\memory[12][3] ),
    .B(_06312_),
    .Y(_07563_)
  );
  NAND _15782_ (
    .A(\memory[27][3] ),
    .B(_06333_),
    .Y(_07564_)
  );
  AND _15783_ (
    .A(_07538_),
    .B(_07549_),
    .Y(_07565_)
  );
  AND _15784_ (
    .A(_07560_),
    .B(_07564_),
    .Y(_07566_)
  );
  AND _15785_ (
    .A(_07531_),
    .B(_07534_),
    .Y(_07567_)
  );
  AND _15786_ (
    .A(_07542_),
    .B(_07563_),
    .Y(_07568_)
  );
  AND _15787_ (
    .A(_07546_),
    .B(_07555_),
    .Y(_07569_)
  );
  AND _15788_ (
    .A(_07540_),
    .B(_07568_),
    .Y(_07570_)
  );
  AND _15789_ (
    .A(_07569_),
    .B(_07570_),
    .Y(_07571_)
  );
  AND _15790_ (
    .A(_07530_),
    .B(_07548_),
    .Y(_07573_)
  );
  AND _15791_ (
    .A(_07553_),
    .B(_07573_),
    .Y(_07574_)
  );
  AND _15792_ (
    .A(_07544_),
    .B(_07557_),
    .Y(_07575_)
  );
  AND _15793_ (
    .A(_07574_),
    .B(_07575_),
    .Y(_07576_)
  );
  AND _15794_ (
    .A(_07571_),
    .B(_07576_),
    .Y(_07577_)
  );
  AND _15795_ (
    .A(_07545_),
    .B(_07558_),
    .Y(_07578_)
  );
  AND _15796_ (
    .A(_07537_),
    .B(_07554_),
    .Y(_07579_)
  );
  AND _15797_ (
    .A(_07533_),
    .B(_07579_),
    .Y(_07580_)
  );
  AND _15798_ (
    .A(_07578_),
    .B(_07580_),
    .Y(_07581_)
  );
  AND _15799_ (
    .A(_07541_),
    .B(_07581_),
    .Y(_07582_)
  );
  AND _15800_ (
    .A(_07552_),
    .B(_07559_),
    .Y(_07584_)
  );
  AND _15801_ (
    .A(_07556_),
    .B(_07584_),
    .Y(_07585_)
  );
  AND _15802_ (
    .A(_07535_),
    .B(_07547_),
    .Y(_07586_)
  );
  AND _15803_ (
    .A(_07567_),
    .B(_07586_),
    .Y(_07587_)
  );
  AND _15804_ (
    .A(_07585_),
    .B(_07587_),
    .Y(_07588_)
  );
  AND _15805_ (
    .A(_07582_),
    .B(_07588_),
    .Y(_07589_)
  );
  AND _15806_ (
    .A(_07543_),
    .B(_07566_),
    .Y(_07590_)
  );
  AND _15807_ (
    .A(_07551_),
    .B(_07590_),
    .Y(_07591_)
  );
  AND _15808_ (
    .A(_07532_),
    .B(_07562_),
    .Y(_07592_)
  );
  AND _15809_ (
    .A(_07536_),
    .B(_07592_),
    .Y(_07593_)
  );
  AND _15810_ (
    .A(_07565_),
    .B(_07593_),
    .Y(_07595_)
  );
  AND _15811_ (
    .A(_07591_),
    .B(_07595_),
    .Y(_07596_)
  );
  AND _15812_ (
    .A(_07589_),
    .B(_07596_),
    .Y(_07597_)
  );
  NAND _15813_ (
    .A(_07577_),
    .B(_07597_),
    .Y(\data_mem_o[27] )
  );
  NAND _15814_ (
    .A(\memory[20][4] ),
    .B(_05754_),
    .Y(_07598_)
  );
  NAND _15815_ (
    .A(\memory[23][4] ),
    .B(_05806_),
    .Y(_07599_)
  );
  NAND _15816_ (
    .A(\memory[15][4] ),
    .B(_06002_),
    .Y(_07600_)
  );
  NAND _15817_ (
    .A(\memory[24][4] ),
    .B(_06023_),
    .Y(_07601_)
  );
  NAND _15818_ (
    .A(\memory[3][4] ),
    .B(_06043_),
    .Y(_07602_)
  );
  NAND _15819_ (
    .A(\memory[8][4] ),
    .B(_05475_),
    .Y(_07603_)
  );
  NAND _15820_ (
    .A(\memory[19][4] ),
    .B(_05558_),
    .Y(_07605_)
  );
  NAND _15821_ (
    .A(\memory[14][4] ),
    .B(_05785_),
    .Y(_07606_)
  );
  NAND _15822_ (
    .A(\memory[7][4] ),
    .B(_05733_),
    .Y(_07607_)
  );
  NAND _15823_ (
    .A(\memory[30][4] ),
    .B(_05847_),
    .Y(_07608_)
  );
  NAND _15824_ (
    .A(\memory[16][4] ),
    .B(_06064_),
    .Y(_07609_)
  );
  NAND _15825_ (
    .A(\memory[12][4] ),
    .B(_06312_),
    .Y(_07610_)
  );
  NAND _15826_ (
    .A(\memory[28][4] ),
    .B(_06291_),
    .Y(_07611_)
  );
  NAND _15827_ (
    .A(\memory[27][4] ),
    .B(_06333_),
    .Y(_07612_)
  );
  NAND _15828_ (
    .A(\memory[29][4] ),
    .B(_05981_),
    .Y(_07613_)
  );
  NAND _15829_ (
    .A(\memory[31][4] ),
    .B(_05826_),
    .Y(_07614_)
  );
  NAND _15830_ (
    .A(\memory[0][4] ),
    .B(_05692_),
    .Y(_07616_)
  );
  AND _15831_ (
    .A(_07614_),
    .B(_07616_),
    .Y(_07617_)
  );
  NAND _15832_ (
    .A(\memory[4][4] ),
    .B(_05599_),
    .Y(_07618_)
  );
  NAND _15833_ (
    .A(\memory[13][4] ),
    .B(_05661_),
    .Y(_07619_)
  );
  NAND _15834_ (
    .A(\memory[10][4] ),
    .B(_06353_),
    .Y(_07620_)
  );
  NAND _15835_ (
    .A(\memory[1][4] ),
    .B(_06188_),
    .Y(_07621_)
  );
  NAND _15836_ (
    .A(\memory[18][4] ),
    .B(_06209_),
    .Y(_07622_)
  );
  NAND _15837_ (
    .A(\memory[2][4] ),
    .B(_06116_),
    .Y(_07623_)
  );
  NAND _15838_ (
    .A(\memory[6][4] ),
    .B(_06147_),
    .Y(_07624_)
  );
  NAND _15839_ (
    .A(\memory[22][4] ),
    .B(_06167_),
    .Y(_07625_)
  );
  NAND _15840_ (
    .A(\memory[26][4] ),
    .B(_06250_),
    .Y(_07627_)
  );
  NAND _15841_ (
    .A(\memory[25][4] ),
    .B(_06395_),
    .Y(_07628_)
  );
  AND _15842_ (
    .A(_07627_),
    .B(_07628_),
    .Y(_07629_)
  );
  NAND _15843_ (
    .A(\memory[9][4] ),
    .B(_06374_),
    .Y(_07630_)
  );
  NAND _15844_ (
    .A(\memory[5][4] ),
    .B(_05961_),
    .Y(_07631_)
  );
  NAND _15845_ (
    .A(\memory[21][4] ),
    .B(_05930_),
    .Y(_07632_)
  );
  NAND _15846_ (
    .A(\memory[11][4] ),
    .B(_05899_),
    .Y(_07633_)
  );
  NAND _15847_ (
    .A(\memory[17][4] ),
    .B(_06085_),
    .Y(_07634_)
  );
  AND _15848_ (
    .A(_07613_),
    .B(_07634_),
    .Y(_07635_)
  );
  AND _15849_ (
    .A(_07624_),
    .B(_07631_),
    .Y(_07636_)
  );
  AND _15850_ (
    .A(_07618_),
    .B(_07636_),
    .Y(_07638_)
  );
  AND _15851_ (
    .A(_07619_),
    .B(_07633_),
    .Y(_07639_)
  );
  AND _15852_ (
    .A(_07612_),
    .B(_07632_),
    .Y(_07640_)
  );
  AND _15853_ (
    .A(_07639_),
    .B(_07640_),
    .Y(_07641_)
  );
  AND _15854_ (
    .A(_07621_),
    .B(_07641_),
    .Y(_07642_)
  );
  AND _15855_ (
    .A(_07606_),
    .B(_07610_),
    .Y(_07643_)
  );
  AND _15856_ (
    .A(_07635_),
    .B(_07643_),
    .Y(_07644_)
  );
  AND _15857_ (
    .A(_07603_),
    .B(_07607_),
    .Y(_07645_)
  );
  AND _15858_ (
    .A(_07623_),
    .B(_07645_),
    .Y(_07646_)
  );
  AND _15859_ (
    .A(_07620_),
    .B(_07646_),
    .Y(_07647_)
  );
  AND _15860_ (
    .A(_07644_),
    .B(_07647_),
    .Y(_07649_)
  );
  AND _15861_ (
    .A(_07642_),
    .B(_07649_),
    .Y(_07650_)
  );
  AND _15862_ (
    .A(_07598_),
    .B(_07601_),
    .Y(_07651_)
  );
  AND _15863_ (
    .A(_07599_),
    .B(_07625_),
    .Y(_07652_)
  );
  AND _15864_ (
    .A(_07608_),
    .B(_07652_),
    .Y(_07653_)
  );
  AND _15865_ (
    .A(_07651_),
    .B(_07653_),
    .Y(_07654_)
  );
  AND _15866_ (
    .A(_07617_),
    .B(_07629_),
    .Y(_07655_)
  );
  AND _15867_ (
    .A(_07654_),
    .B(_07655_),
    .Y(_07656_)
  );
  AND _15868_ (
    .A(_07605_),
    .B(_07611_),
    .Y(_07657_)
  );
  AND _15869_ (
    .A(_07622_),
    .B(_07657_),
    .Y(_07658_)
  );
  AND _15870_ (
    .A(_07600_),
    .B(_07609_),
    .Y(_07660_)
  );
  AND _15871_ (
    .A(_07602_),
    .B(_07630_),
    .Y(_07661_)
  );
  AND _15872_ (
    .A(_07660_),
    .B(_07661_),
    .Y(_07662_)
  );
  AND _15873_ (
    .A(_07658_),
    .B(_07662_),
    .Y(_07663_)
  );
  AND _15874_ (
    .A(_07656_),
    .B(_07663_),
    .Y(_07664_)
  );
  AND _15875_ (
    .A(_07650_),
    .B(_07664_),
    .Y(_07665_)
  );
  NAND _15876_ (
    .A(_07638_),
    .B(_07665_),
    .Y(\data_mem_o[28] )
  );
  NAND _15877_ (
    .A(\memory[30][5] ),
    .B(_05847_),
    .Y(_07666_)
  );
  NAND _15878_ (
    .A(\memory[14][5] ),
    .B(_05785_),
    .Y(_07667_)
  );
  NAND _15879_ (
    .A(\memory[7][5] ),
    .B(_05733_),
    .Y(_07668_)
  );
  NAND _15880_ (
    .A(\memory[19][5] ),
    .B(_05558_),
    .Y(_07670_)
  );
  NAND _15881_ (
    .A(\memory[15][5] ),
    .B(_06002_),
    .Y(_07671_)
  );
  NAND _15882_ (
    .A(\memory[13][5] ),
    .B(_05661_),
    .Y(_07672_)
  );
  NAND _15883_ (
    .A(\memory[23][5] ),
    .B(_05806_),
    .Y(_07673_)
  );
  NAND _15884_ (
    .A(\memory[24][5] ),
    .B(_06023_),
    .Y(_07674_)
  );
  NAND _15885_ (
    .A(\memory[3][5] ),
    .B(_06043_),
    .Y(_07675_)
  );
  NAND _15886_ (
    .A(\memory[8][5] ),
    .B(_05475_),
    .Y(_07676_)
  );
  NAND _15887_ (
    .A(\memory[16][5] ),
    .B(_06064_),
    .Y(_07677_)
  );
  NAND _15888_ (
    .A(\memory[12][5] ),
    .B(_06312_),
    .Y(_07678_)
  );
  NAND _15889_ (
    .A(\memory[10][5] ),
    .B(_06353_),
    .Y(_07679_)
  );
  NAND _15890_ (
    .A(\memory[27][5] ),
    .B(_06333_),
    .Y(_07681_)
  );
  NAND _15891_ (
    .A(\memory[29][5] ),
    .B(_05981_),
    .Y(_07682_)
  );
  NAND _15892_ (
    .A(\memory[31][5] ),
    .B(_05826_),
    .Y(_07683_)
  );
  NAND _15893_ (
    .A(\memory[0][5] ),
    .B(_05692_),
    .Y(_07684_)
  );
  AND _15894_ (
    .A(_07683_),
    .B(_07684_),
    .Y(_07685_)
  );
  NAND _15895_ (
    .A(\memory[4][5] ),
    .B(_05599_),
    .Y(_07686_)
  );
  NAND _15896_ (
    .A(\memory[20][5] ),
    .B(_05754_),
    .Y(_07687_)
  );
  NAND _15897_ (
    .A(\memory[28][5] ),
    .B(_06291_),
    .Y(_07688_)
  );
  NAND _15898_ (
    .A(\memory[1][5] ),
    .B(_06188_),
    .Y(_07689_)
  );
  NAND _15899_ (
    .A(\memory[6][5] ),
    .B(_06147_),
    .Y(_07690_)
  );
  NAND _15900_ (
    .A(\memory[22][5] ),
    .B(_06167_),
    .Y(_07692_)
  );
  NAND _15901_ (
    .A(\memory[2][5] ),
    .B(_06116_),
    .Y(_07693_)
  );
  NAND _15902_ (
    .A(\memory[18][5] ),
    .B(_06209_),
    .Y(_07694_)
  );
  NAND _15903_ (
    .A(\memory[21][5] ),
    .B(_05930_),
    .Y(_07695_)
  );
  NAND _15904_ (
    .A(\memory[25][5] ),
    .B(_06395_),
    .Y(_07696_)
  );
  NAND _15905_ (
    .A(\memory[9][5] ),
    .B(_06374_),
    .Y(_07697_)
  );
  NAND _15906_ (
    .A(\memory[5][5] ),
    .B(_05961_),
    .Y(_07698_)
  );
  NAND _15907_ (
    .A(\memory[11][5] ),
    .B(_05899_),
    .Y(_07699_)
  );
  NAND _15908_ (
    .A(\memory[17][5] ),
    .B(_06085_),
    .Y(_07700_)
  );
  NAND _15909_ (
    .A(\memory[26][5] ),
    .B(_06250_),
    .Y(_07701_)
  );
  AND _15910_ (
    .A(_07696_),
    .B(_07701_),
    .Y(_07703_)
  );
  AND _15911_ (
    .A(_07682_),
    .B(_07700_),
    .Y(_07704_)
  );
  AND _15912_ (
    .A(_07690_),
    .B(_07698_),
    .Y(_07705_)
  );
  AND _15913_ (
    .A(_07686_),
    .B(_07705_),
    .Y(_07706_)
  );
  AND _15914_ (
    .A(_07672_),
    .B(_07699_),
    .Y(_07707_)
  );
  AND _15915_ (
    .A(_07681_),
    .B(_07695_),
    .Y(_07708_)
  );
  AND _15916_ (
    .A(_07707_),
    .B(_07708_),
    .Y(_07709_)
  );
  AND _15917_ (
    .A(_07689_),
    .B(_07709_),
    .Y(_07710_)
  );
  AND _15918_ (
    .A(_07667_),
    .B(_07678_),
    .Y(_07711_)
  );
  AND _15919_ (
    .A(_07704_),
    .B(_07711_),
    .Y(_07712_)
  );
  AND _15920_ (
    .A(_07668_),
    .B(_07676_),
    .Y(_07714_)
  );
  AND _15921_ (
    .A(_07693_),
    .B(_07714_),
    .Y(_07715_)
  );
  AND _15922_ (
    .A(_07679_),
    .B(_07715_),
    .Y(_07716_)
  );
  AND _15923_ (
    .A(_07712_),
    .B(_07716_),
    .Y(_07717_)
  );
  AND _15924_ (
    .A(_07710_),
    .B(_07717_),
    .Y(_07718_)
  );
  AND _15925_ (
    .A(_07674_),
    .B(_07687_),
    .Y(_07719_)
  );
  AND _15926_ (
    .A(_07673_),
    .B(_07692_),
    .Y(_07720_)
  );
  AND _15927_ (
    .A(_07666_),
    .B(_07720_),
    .Y(_07721_)
  );
  AND _15928_ (
    .A(_07719_),
    .B(_07721_),
    .Y(_07722_)
  );
  AND _15929_ (
    .A(_07685_),
    .B(_07703_),
    .Y(_07723_)
  );
  AND _15930_ (
    .A(_07722_),
    .B(_07723_),
    .Y(_07725_)
  );
  AND _15931_ (
    .A(_07670_),
    .B(_07688_),
    .Y(_07726_)
  );
  AND _15932_ (
    .A(_07694_),
    .B(_07726_),
    .Y(_07727_)
  );
  AND _15933_ (
    .A(_07671_),
    .B(_07677_),
    .Y(_07728_)
  );
  AND _15934_ (
    .A(_07675_),
    .B(_07697_),
    .Y(_07729_)
  );
  AND _15935_ (
    .A(_07728_),
    .B(_07729_),
    .Y(_07730_)
  );
  AND _15936_ (
    .A(_07727_),
    .B(_07730_),
    .Y(_07731_)
  );
  AND _15937_ (
    .A(_07725_),
    .B(_07731_),
    .Y(_07732_)
  );
  AND _15938_ (
    .A(_07718_),
    .B(_07732_),
    .Y(_07733_)
  );
  NAND _15939_ (
    .A(_07706_),
    .B(_07733_),
    .Y(\data_mem_o[29] )
  );
  NAND _15940_ (
    .A(\memory[14][6] ),
    .B(_05785_),
    .Y(_07735_)
  );
  NAND _15941_ (
    .A(\memory[8][6] ),
    .B(_05475_),
    .Y(_07736_)
  );
  NAND _15942_ (
    .A(\memory[4][6] ),
    .B(_05599_),
    .Y(_07737_)
  );
  NAND _15943_ (
    .A(\memory[20][6] ),
    .B(_05754_),
    .Y(_07738_)
  );
  NAND _15944_ (
    .A(\memory[0][6] ),
    .B(_05692_),
    .Y(_07739_)
  );
  NAND _15945_ (
    .A(\memory[24][6] ),
    .B(_06023_),
    .Y(_07740_)
  );
  NAND _15946_ (
    .A(\memory[19][6] ),
    .B(_05558_),
    .Y(_07741_)
  );
  NAND _15947_ (
    .A(\memory[23][6] ),
    .B(_05806_),
    .Y(_07742_)
  );
  NAND _15948_ (
    .A(\memory[15][6] ),
    .B(_06002_),
    .Y(_07743_)
  );
  NAND _15949_ (
    .A(\memory[7][6] ),
    .B(_05733_),
    .Y(_07744_)
  );
  NAND _15950_ (
    .A(\memory[31][6] ),
    .B(_05826_),
    .Y(_07746_)
  );
  NAND _15951_ (
    .A(\memory[26][6] ),
    .B(_06250_),
    .Y(_07747_)
  );
  NAND _15952_ (
    .A(\memory[25][6] ),
    .B(_06395_),
    .Y(_07748_)
  );
  AND _15953_ (
    .A(_07747_),
    .B(_07748_),
    .Y(_07749_)
  );
  NAND _15954_ (
    .A(\memory[28][6] ),
    .B(_06291_),
    .Y(_07750_)
  );
  NAND _15955_ (
    .A(\memory[21][6] ),
    .B(_05930_),
    .Y(_07751_)
  );
  NAND _15956_ (
    .A(\memory[30][6] ),
    .B(_05847_),
    .Y(_07752_)
  );
  NAND _15957_ (
    .A(\memory[16][6] ),
    .B(_06064_),
    .Y(_07753_)
  );
  NAND _15958_ (
    .A(\memory[3][6] ),
    .B(_06043_),
    .Y(_07754_)
  );
  NAND _15959_ (
    .A(\memory[13][6] ),
    .B(_05661_),
    .Y(_07755_)
  );
  NAND _15960_ (
    .A(\memory[17][6] ),
    .B(_06085_),
    .Y(_07757_)
  );
  NAND _15961_ (
    .A(\memory[2][6] ),
    .B(_06116_),
    .Y(_07758_)
  );
  NAND _15962_ (
    .A(\memory[22][6] ),
    .B(_06167_),
    .Y(_07759_)
  );
  NAND _15963_ (
    .A(\memory[6][6] ),
    .B(_06147_),
    .Y(_07760_)
  );
  NAND _15964_ (
    .A(\memory[1][6] ),
    .B(_06188_),
    .Y(_07761_)
  );
  NAND _15965_ (
    .A(\memory[18][6] ),
    .B(_06209_),
    .Y(_07762_)
  );
  NAND _15966_ (
    .A(\memory[10][6] ),
    .B(_06353_),
    .Y(_07763_)
  );
  NAND _15967_ (
    .A(\memory[9][6] ),
    .B(_06374_),
    .Y(_07764_)
  );
  NAND _15968_ (
    .A(\memory[29][6] ),
    .B(_05981_),
    .Y(_07765_)
  );
  NAND _15969_ (
    .A(\memory[12][6] ),
    .B(_06312_),
    .Y(_07766_)
  );
  NAND _15970_ (
    .A(\memory[27][6] ),
    .B(_06333_),
    .Y(_07768_)
  );
  NAND _15971_ (
    .A(\memory[5][6] ),
    .B(_05961_),
    .Y(_07769_)
  );
  NAND _15972_ (
    .A(\memory[11][6] ),
    .B(_05899_),
    .Y(_07770_)
  );
  AND _15973_ (
    .A(_07743_),
    .B(_07753_),
    .Y(_07771_)
  );
  AND _15974_ (
    .A(_07736_),
    .B(_07744_),
    .Y(_07772_)
  );
  AND _15975_ (
    .A(_07751_),
    .B(_07765_),
    .Y(_07773_)
  );
  AND _15976_ (
    .A(_07735_),
    .B(_07766_),
    .Y(_07774_)
  );
  AND _15977_ (
    .A(_07757_),
    .B(_07774_),
    .Y(_07775_)
  );
  AND _15978_ (
    .A(_07758_),
    .B(_07772_),
    .Y(_07776_)
  );
  AND _15979_ (
    .A(_07763_),
    .B(_07776_),
    .Y(_07777_)
  );
  AND _15980_ (
    .A(_07761_),
    .B(_07777_),
    .Y(_07779_)
  );
  AND _15981_ (
    .A(_07775_),
    .B(_07779_),
    .Y(_07780_)
  );
  AND _15982_ (
    .A(_07738_),
    .B(_07740_),
    .Y(_07781_)
  );
  AND _15983_ (
    .A(_07742_),
    .B(_07759_),
    .Y(_07782_)
  );
  AND _15984_ (
    .A(_07752_),
    .B(_07782_),
    .Y(_07783_)
  );
  AND _15985_ (
    .A(_07781_),
    .B(_07783_),
    .Y(_07784_)
  );
  AND _15986_ (
    .A(_07739_),
    .B(_07746_),
    .Y(_07785_)
  );
  AND _15987_ (
    .A(_07749_),
    .B(_07785_),
    .Y(_07786_)
  );
  AND _15988_ (
    .A(_07784_),
    .B(_07786_),
    .Y(_07787_)
  );
  AND _15989_ (
    .A(_07741_),
    .B(_07750_),
    .Y(_07788_)
  );
  AND _15990_ (
    .A(_07762_),
    .B(_07788_),
    .Y(_07790_)
  );
  AND _15991_ (
    .A(_07754_),
    .B(_07764_),
    .Y(_07791_)
  );
  AND _15992_ (
    .A(_07771_),
    .B(_07791_),
    .Y(_07792_)
  );
  AND _15993_ (
    .A(_07790_),
    .B(_07792_),
    .Y(_07793_)
  );
  AND _15994_ (
    .A(_07787_),
    .B(_07793_),
    .Y(_07794_)
  );
  AND _15995_ (
    .A(_07780_),
    .B(_07794_),
    .Y(_07795_)
  );
  AND _15996_ (
    .A(_07760_),
    .B(_07769_),
    .Y(_07796_)
  );
  AND _15997_ (
    .A(_07737_),
    .B(_07796_),
    .Y(_07797_)
  );
  AND _15998_ (
    .A(_07755_),
    .B(_07770_),
    .Y(_07798_)
  );
  AND _15999_ (
    .A(_07768_),
    .B(_07773_),
    .Y(_07799_)
  );
  AND _16000_ (
    .A(_07798_),
    .B(_07799_),
    .Y(_07801_)
  );
  AND _16001_ (
    .A(_07797_),
    .B(_07801_),
    .Y(_07802_)
  );
  NAND _16002_ (
    .A(_07795_),
    .B(_07802_),
    .Y(\data_mem_o[30] )
  );
  NAND _16003_ (
    .A(\memory[14][7] ),
    .B(_05785_),
    .Y(_07803_)
  );
  NAND _16004_ (
    .A(\memory[8][7] ),
    .B(_05475_),
    .Y(_07804_)
  );
  NAND _16005_ (
    .A(\memory[4][7] ),
    .B(_05599_),
    .Y(_07805_)
  );
  NAND _16006_ (
    .A(\memory[20][7] ),
    .B(_05754_),
    .Y(_07806_)
  );
  NAND _16007_ (
    .A(\memory[0][7] ),
    .B(_05692_),
    .Y(_07807_)
  );
  NAND _16008_ (
    .A(\memory[24][7] ),
    .B(_06023_),
    .Y(_07808_)
  );
  NAND _16009_ (
    .A(\memory[19][7] ),
    .B(_05558_),
    .Y(_07809_)
  );
  NAND _16010_ (
    .A(\memory[23][7] ),
    .B(_05806_),
    .Y(_07811_)
  );
  NAND _16011_ (
    .A(\memory[15][7] ),
    .B(_06002_),
    .Y(_07812_)
  );
  NAND _16012_ (
    .A(\memory[7][7] ),
    .B(_05733_),
    .Y(_07813_)
  );
  NAND _16013_ (
    .A(\memory[31][7] ),
    .B(_05826_),
    .Y(_07814_)
  );
  NAND _16014_ (
    .A(\memory[26][7] ),
    .B(_06250_),
    .Y(_07815_)
  );
  NAND _16015_ (
    .A(\memory[25][7] ),
    .B(_06395_),
    .Y(_07816_)
  );
  AND _16016_ (
    .A(_07815_),
    .B(_07816_),
    .Y(_07817_)
  );
  NAND _16017_ (
    .A(\memory[28][7] ),
    .B(_06291_),
    .Y(_07818_)
  );
  NAND _16018_ (
    .A(\memory[21][7] ),
    .B(_05930_),
    .Y(_07819_)
  );
  NAND _16019_ (
    .A(\memory[30][7] ),
    .B(_05847_),
    .Y(_07820_)
  );
  NAND _16020_ (
    .A(\memory[16][7] ),
    .B(_06064_),
    .Y(_07822_)
  );
  NAND _16021_ (
    .A(\memory[3][7] ),
    .B(_06043_),
    .Y(_07823_)
  );
  NAND _16022_ (
    .A(\memory[13][7] ),
    .B(_05661_),
    .Y(_07824_)
  );
  NAND _16023_ (
    .A(\memory[17][7] ),
    .B(_06085_),
    .Y(_07825_)
  );
  NAND _16024_ (
    .A(\memory[2][7] ),
    .B(_06116_),
    .Y(_07826_)
  );
  NAND _16025_ (
    .A(\memory[22][7] ),
    .B(_06167_),
    .Y(_07827_)
  );
  NAND _16026_ (
    .A(\memory[6][7] ),
    .B(_06147_),
    .Y(_07828_)
  );
  NAND _16027_ (
    .A(\memory[1][7] ),
    .B(_06188_),
    .Y(_07829_)
  );
  NAND _16028_ (
    .A(\memory[18][7] ),
    .B(_06209_),
    .Y(_07830_)
  );
  NAND _16029_ (
    .A(\memory[10][7] ),
    .B(_06353_),
    .Y(_07831_)
  );
  NAND _16030_ (
    .A(\memory[9][7] ),
    .B(_06374_),
    .Y(_07833_)
  );
  NAND _16031_ (
    .A(\memory[29][7] ),
    .B(_05981_),
    .Y(_07834_)
  );
  NAND _16032_ (
    .A(\memory[12][7] ),
    .B(_06312_),
    .Y(_07835_)
  );
  NAND _16033_ (
    .A(\memory[27][7] ),
    .B(_06333_),
    .Y(_07836_)
  );
  NAND _16034_ (
    .A(\memory[5][7] ),
    .B(_05961_),
    .Y(_07837_)
  );
  NAND _16035_ (
    .A(\memory[11][7] ),
    .B(_05899_),
    .Y(_07838_)
  );
  AND _16036_ (
    .A(_07812_),
    .B(_07822_),
    .Y(_07839_)
  );
  AND _16037_ (
    .A(_07804_),
    .B(_07813_),
    .Y(_07840_)
  );
  AND _16038_ (
    .A(_07819_),
    .B(_07834_),
    .Y(_07841_)
  );
  AND _16039_ (
    .A(_07803_),
    .B(_07835_),
    .Y(_07842_)
  );
  AND _16040_ (
    .A(_07825_),
    .B(_07842_),
    .Y(_07844_)
  );
  AND _16041_ (
    .A(_07826_),
    .B(_07840_),
    .Y(_07845_)
  );
  AND _16042_ (
    .A(_07831_),
    .B(_07845_),
    .Y(_07846_)
  );
  AND _16043_ (
    .A(_07829_),
    .B(_07846_),
    .Y(_07847_)
  );
  AND _16044_ (
    .A(_07844_),
    .B(_07847_),
    .Y(_07848_)
  );
  AND _16045_ (
    .A(_07806_),
    .B(_07808_),
    .Y(_07849_)
  );
  AND _16046_ (
    .A(_07811_),
    .B(_07827_),
    .Y(_07850_)
  );
  AND _16047_ (
    .A(_07820_),
    .B(_07850_),
    .Y(_07851_)
  );
  AND _16048_ (
    .A(_07849_),
    .B(_07851_),
    .Y(_07852_)
  );
  AND _16049_ (
    .A(_07807_),
    .B(_07814_),
    .Y(_07853_)
  );
  AND _16050_ (
    .A(_07817_),
    .B(_07853_),
    .Y(_07855_)
  );
  AND _16051_ (
    .A(_07852_),
    .B(_07855_),
    .Y(_07856_)
  );
  AND _16052_ (
    .A(_07809_),
    .B(_07818_),
    .Y(_07857_)
  );
  AND _16053_ (
    .A(_07830_),
    .B(_07857_),
    .Y(_07858_)
  );
  AND _16054_ (
    .A(_07823_),
    .B(_07833_),
    .Y(_07859_)
  );
  AND _16055_ (
    .A(_07839_),
    .B(_07859_),
    .Y(_07860_)
  );
  AND _16056_ (
    .A(_07858_),
    .B(_07860_),
    .Y(_07861_)
  );
  AND _16057_ (
    .A(_07856_),
    .B(_07861_),
    .Y(_07862_)
  );
  AND _16058_ (
    .A(_07848_),
    .B(_07862_),
    .Y(_07863_)
  );
  AND _16059_ (
    .A(_07828_),
    .B(_07837_),
    .Y(_07864_)
  );
  AND _16060_ (
    .A(_07805_),
    .B(_07864_),
    .Y(_07866_)
  );
  AND _16061_ (
    .A(_07824_),
    .B(_07838_),
    .Y(_07867_)
  );
  AND _16062_ (
    .A(_07836_),
    .B(_07841_),
    .Y(_07868_)
  );
  AND _16063_ (
    .A(_07867_),
    .B(_07868_),
    .Y(_07869_)
  );
  AND _16064_ (
    .A(_07866_),
    .B(_07869_),
    .Y(_07870_)
  );
  NAND _16065_ (
    .A(_07863_),
    .B(_07870_),
    .Y(\data_mem_o[31] )
  );
endmodule

module EX_Mem (
MemRead_i, 
MemRead_o, 
MemToReg_i, 
MemToReg_o, 
MemWrite_i, 
MemWrite_o, 
RegWrite_i, 
RegWrite_o, 
\ALUResult_i[0], 
\ALUResult_i[10], 
\ALUResult_i[11], 
\ALUResult_i[12], 
\ALUResult_i[13], 
\ALUResult_i[14], 
\ALUResult_i[15], 
\ALUResult_i[16], 
\ALUResult_i[17], 
\ALUResult_i[18], 
\ALUResult_i[19], 
\ALUResult_i[1], 
\ALUResult_i[20], 
\ALUResult_i[21], 
\ALUResult_i[22], 
\ALUResult_i[23], 
\ALUResult_i[24], 
\ALUResult_i[25], 
\ALUResult_i[26], 
\ALUResult_i[27], 
\ALUResult_i[28], 
\ALUResult_i[29], 
\ALUResult_i[2], 
\ALUResult_i[30], 
\ALUResult_i[31], 
\ALUResult_i[3], 
\ALUResult_i[4], 
\ALUResult_i[5], 
\ALUResult_i[6], 
\ALUResult_i[7], 
\ALUResult_i[8], 
\ALUResult_i[9], 
\ALUResult_o[0], 
\ALUResult_o[10], 
\ALUResult_o[11], 
\ALUResult_o[12], 
\ALUResult_o[13], 
\ALUResult_o[14], 
\ALUResult_o[15], 
\ALUResult_o[16], 
\ALUResult_o[17], 
\ALUResult_o[18], 
\ALUResult_o[19], 
\ALUResult_o[1], 
\ALUResult_o[20], 
\ALUResult_o[21], 
\ALUResult_o[22], 
\ALUResult_o[23], 
\ALUResult_o[24], 
\ALUResult_o[25], 
\ALUResult_o[26], 
\ALUResult_o[27], 
\ALUResult_o[28], 
\ALUResult_o[29], 
\ALUResult_o[2], 
\ALUResult_o[30], 
\ALUResult_o[31], 
\ALUResult_o[3], 
\ALUResult_o[4], 
\ALUResult_o[5], 
\ALUResult_o[6], 
\ALUResult_o[7], 
\ALUResult_o[8], 
\ALUResult_o[9], 
\RDData_i[0], 
\RDData_i[10], 
\RDData_i[11], 
\RDData_i[12], 
\RDData_i[13], 
\RDData_i[14], 
\RDData_i[15], 
\RDData_i[16], 
\RDData_i[17], 
\RDData_i[18], 
\RDData_i[19], 
\RDData_i[1], 
\RDData_i[20], 
\RDData_i[21], 
\RDData_i[22], 
\RDData_i[23], 
\RDData_i[24], 
\RDData_i[25], 
\RDData_i[26], 
\RDData_i[27], 
\RDData_i[28], 
\RDData_i[29], 
\RDData_i[2], 
\RDData_i[30], 
\RDData_i[31], 
\RDData_i[3], 
\RDData_i[4], 
\RDData_i[5], 
\RDData_i[6], 
\RDData_i[7], 
\RDData_i[8], 
\RDData_i[9], 
\RDData_o[0], 
\RDData_o[10], 
\RDData_o[11], 
\RDData_o[12], 
\RDData_o[13], 
\RDData_o[14], 
\RDData_o[15], 
\RDData_o[16], 
\RDData_o[17], 
\RDData_o[18], 
\RDData_o[19], 
\RDData_o[1], 
\RDData_o[20], 
\RDData_o[21], 
\RDData_o[22], 
\RDData_o[23], 
\RDData_o[24], 
\RDData_o[25], 
\RDData_o[26], 
\RDData_o[27], 
\RDData_o[28], 
\RDData_o[29], 
\RDData_o[2], 
\RDData_o[30], 
\RDData_o[31], 
\RDData_o[3], 
\RDData_o[4], 
\RDData_o[5], 
\RDData_o[6], 
\RDData_o[7], 
\RDData_o[8], 
\RDData_o[9], 
\RDaddr_i[0], 
\RDaddr_i[1], 
\RDaddr_i[2], 
\RDaddr_i[3], 
\RDaddr_i[4], 
\RDaddr_o[0], 
\RDaddr_o[1], 
\RDaddr_o[2], 
\RDaddr_o[3], 
\RDaddr_o[4], 
\VALUResult_i[0], 
\VALUResult_i[10], 
\VALUResult_i[11], 
\VALUResult_i[12], 
\VALUResult_i[13], 
\VALUResult_i[14], 
\VALUResult_i[15], 
\VALUResult_i[16], 
\VALUResult_i[17], 
\VALUResult_i[18], 
\VALUResult_i[19], 
\VALUResult_i[1], 
\VALUResult_i[20], 
\VALUResult_i[21], 
\VALUResult_i[22], 
\VALUResult_i[23], 
\VALUResult_i[24], 
\VALUResult_i[25], 
\VALUResult_i[26], 
\VALUResult_i[27], 
\VALUResult_i[28], 
\VALUResult_i[29], 
\VALUResult_i[2], 
\VALUResult_i[30], 
\VALUResult_i[31], 
\VALUResult_i[3], 
\VALUResult_i[4], 
\VALUResult_i[5], 
\VALUResult_i[6], 
\VALUResult_i[7], 
\VALUResult_i[8], 
\VALUResult_i[9], 
\VALUResult_o[0], 
\VALUResult_o[10], 
\VALUResult_o[11], 
\VALUResult_o[12], 
\VALUResult_o[13], 
\VALUResult_o[14], 
\VALUResult_o[15], 
\VALUResult_o[16], 
\VALUResult_o[17], 
\VALUResult_o[18], 
\VALUResult_o[19], 
\VALUResult_o[1], 
\VALUResult_o[20], 
\VALUResult_o[21], 
\VALUResult_o[22], 
\VALUResult_o[23], 
\VALUResult_o[24], 
\VALUResult_o[25], 
\VALUResult_o[26], 
\VALUResult_o[27], 
\VALUResult_o[28], 
\VALUResult_o[29], 
\VALUResult_o[2], 
\VALUResult_o[30], 
\VALUResult_o[31], 
\VALUResult_o[3], 
\VALUResult_o[4], 
\VALUResult_o[5], 
\VALUResult_o[6], 
\VALUResult_o[7], 
\VALUResult_o[8], 
\VALUResult_o[9], 
\instr_i[0], 
\instr_i[10], 
\instr_i[11], 
\instr_i[12], 
\instr_i[13], 
\instr_i[14], 
\instr_i[15], 
\instr_i[16], 
\instr_i[17], 
\instr_i[18], 
\instr_i[19], 
\instr_i[1], 
\instr_i[20], 
\instr_i[21], 
\instr_i[22], 
\instr_i[23], 
\instr_i[24], 
\instr_i[25], 
\instr_i[26], 
\instr_i[27], 
\instr_i[28], 
\instr_i[29], 
\instr_i[2], 
\instr_i[30], 
\instr_i[31], 
\instr_i[3], 
\instr_i[4], 
\instr_i[5], 
\instr_i[6], 
\instr_i[7], 
\instr_i[8], 
\instr_i[9], 
\instr_o[0], 
\instr_o[10], 
\instr_o[11], 
\instr_o[12], 
\instr_o[13], 
\instr_o[14], 
\instr_o[15], 
\instr_o[16], 
\instr_o[17], 
\instr_o[18], 
\instr_o[19], 
\instr_o[1], 
\instr_o[20], 
\instr_o[21], 
\instr_o[22], 
\instr_o[23], 
\instr_o[24], 
\instr_o[25], 
\instr_o[26], 
\instr_o[27], 
\instr_o[28], 
\instr_o[29], 
\instr_o[2], 
\instr_o[30], 
\instr_o[31], 
\instr_o[3], 
\instr_o[4], 
\instr_o[5], 
\instr_o[6], 
\instr_o[7], 
\instr_o[8], 
\instr_o[9], 
\pc_i[0], 
\pc_i[10], 
\pc_i[11], 
\pc_i[12], 
\pc_i[13], 
\pc_i[14], 
\pc_i[15], 
\pc_i[16], 
\pc_i[17], 
\pc_i[18], 
\pc_i[19], 
\pc_i[1], 
\pc_i[20], 
\pc_i[21], 
\pc_i[22], 
\pc_i[23], 
\pc_i[24], 
\pc_i[25], 
\pc_i[26], 
\pc_i[27], 
\pc_i[28], 
\pc_i[29], 
\pc_i[2], 
\pc_i[30], 
\pc_i[31], 
\pc_i[3], 
\pc_i[4], 
\pc_i[5], 
\pc_i[6], 
\pc_i[7], 
\pc_i[8], 
\pc_i[9], 
\pc_o[0], 
\pc_o[10], 
\pc_o[11], 
\pc_o[12], 
\pc_o[13], 
\pc_o[14], 
\pc_o[15], 
\pc_o[16], 
\pc_o[17], 
\pc_o[18], 
\pc_o[19], 
\pc_o[1], 
\pc_o[20], 
\pc_o[21], 
\pc_o[22], 
\pc_o[23], 
\pc_o[24], 
\pc_o[25], 
\pc_o[26], 
\pc_o[27], 
\pc_o[28], 
\pc_o[29], 
\pc_o[2], 
\pc_o[30], 
\pc_o[31], 
\pc_o[3], 
\pc_o[4], 
\pc_o[5], 
\pc_o[6], 
\pc_o[7], 
\pc_o[8], 
\pc_o[9], 
clk_i, 
start_i, 
zero_i, 
zero_o,
);
  wire _000_ ;
  wire _001_ ;
  wire _002_ ;
  wire _003_ ;
  wire _004_ ;
  wire _005_ ;
  wire _006_ ;
  wire _007_ ;
  wire _008_ ;
  wire _009_ ;
  wire _010_ ;
  wire _011_ ;
  wire _012_ ;
  wire _013_ ;
  wire _014_ ;
  wire _015_ ;
  wire _016_ ;
  wire _017_ ;
  wire _018_ ;
  wire _019_ ;
  wire _020_ ;
  wire _021_ ;
  wire _022_ ;
  wire _023_ ;
  wire _024_ ;
  wire _025_ ;
  wire _026_ ;
  wire _027_ ;
  wire _028_ ;
  wire _029_ ;
  wire _030_ ;
  wire _031_ ;
  wire _032_ ;
  wire _033_ ;
  wire _034_ ;
  wire _035_ ;
  wire _036_ ;
  wire _037_ ;
  wire _038_ ;
  wire _039_ ;
  wire _040_ ;
  wire _041_ ;
  wire _042_ ;
  wire _043_ ;
  wire _044_ ;
  wire _045_ ;
  wire _046_ ;
  wire _047_ ;
  wire _048_ ;
  wire _049_ ;
  wire _050_ ;
  wire _051_ ;
  wire _052_ ;
  wire _053_ ;
  wire _054_ ;
  wire _055_ ;
  wire _056_ ;
  wire _057_ ;
  wire _058_ ;
  wire _059_ ;
  wire _060_ ;
  wire _061_ ;
  wire _062_ ;
  wire _063_ ;
  wire _064_ ;
  wire _065_ ;
  wire _066_ ;
  wire _067_ ;
  wire _068_ ;
  wire _069_ ;
  wire _070_ ;
  wire _071_ ;
  wire _072_ ;
  wire _073_ ;
  wire _074_ ;
  wire _075_ ;
  wire _076_ ;
  wire _077_ ;
  wire _078_ ;
  wire _079_ ;
  wire _080_ ;
  wire _081_ ;
  wire _082_ ;
  wire _083_ ;
  wire _084_ ;
  wire _085_ ;
  wire _086_ ;
  wire _087_ ;
  wire _088_ ;
  wire _089_ ;
  wire _090_ ;
  wire _091_ ;
  wire _092_ ;
  wire _093_ ;
  wire _094_ ;
  wire _095_ ;
  wire _096_ ;
  wire _097_ ;
  wire _098_ ;
  wire _099_ ;
  wire _100_ ;
  wire _101_ ;
  wire _102_ ;
  wire _103_ ;
  wire _104_ ;
  wire _105_ ;
  wire _106_ ;
  wire _107_ ;
  wire _108_ ;
  wire _109_ ;
  wire _110_ ;
  wire _111_ ;
  wire _112_ ;
  wire _113_ ;
  wire _114_ ;
  wire _115_ ;
  wire _116_ ;
  wire _117_ ;
  wire _118_ ;
  wire _119_ ;
  wire _120_ ;
  wire _121_ ;
  wire _122_ ;
  wire _123_ ;
  wire _124_ ;
  wire _125_ ;
  wire _126_ ;
  wire _127_ ;
  wire _128_ ;
  wire _129_ ;
  wire _130_ ;
  wire _131_ ;
  wire _132_ ;
  wire _133_ ;
  wire _134_ ;
  wire _135_ ;
  wire _136_ ;
  wire _137_ ;
  wire _138_ ;
  wire _139_ ;
  wire _140_ ;
  wire _141_ ;
  wire _142_ ;
  wire _143_ ;
  wire _144_ ;
  wire _145_ ;
  wire _146_ ;
  wire _147_ ;
  wire _148_ ;
  wire _149_ ;
  wire _150_ ;
  wire _151_ ;
  wire _152_ ;
  wire _153_ ;
  wire _154_ ;
  wire _155_ ;
  wire _156_ ;
  wire _157_ ;
  wire _158_ ;
  wire _159_ ;
  wire _160_ ;
  wire _161_ ;
  wire _162_ ;
  wire _163_ ;
  wire _164_ ;
  wire _165_ ;
  wire _166_ ;
  wire _167_ ;
  wire _168_ ;
  wire _169_ ;
  input MemRead_i ;
  input MemRead_o ;
  input MemToReg_i ;
  input MemToReg_o ;
  input MemWrite_i ;
  input MemWrite_o ;
  input RegWrite_i ;
  input RegWrite_o ;
  input \ALUResult_i[0] ;
  input \ALUResult_i[10] ;
  input \ALUResult_i[11] ;
  input \ALUResult_i[12] ;
  input \ALUResult_i[13] ;
  input \ALUResult_i[14] ;
  input \ALUResult_i[15] ;
  input \ALUResult_i[16] ;
  input \ALUResult_i[17] ;
  input \ALUResult_i[18] ;
  input \ALUResult_i[19] ;
  input \ALUResult_i[1] ;
  input \ALUResult_i[20] ;
  input \ALUResult_i[21] ;
  input \ALUResult_i[22] ;
  input \ALUResult_i[23] ;
  input \ALUResult_i[24] ;
  input \ALUResult_i[25] ;
  input \ALUResult_i[26] ;
  input \ALUResult_i[27] ;
  input \ALUResult_i[28] ;
  input \ALUResult_i[29] ;
  input \ALUResult_i[2] ;
  input \ALUResult_i[30] ;
  input \ALUResult_i[31] ;
  input \ALUResult_i[3] ;
  input \ALUResult_i[4] ;
  input \ALUResult_i[5] ;
  input \ALUResult_i[6] ;
  input \ALUResult_i[7] ;
  input \ALUResult_i[8] ;
  input \ALUResult_i[9] ;
  input \ALUResult_o[0] ;
  input \ALUResult_o[10] ;
  input \ALUResult_o[11] ;
  input \ALUResult_o[12] ;
  input \ALUResult_o[13] ;
  input \ALUResult_o[14] ;
  input \ALUResult_o[15] ;
  input \ALUResult_o[16] ;
  input \ALUResult_o[17] ;
  input \ALUResult_o[18] ;
  input \ALUResult_o[19] ;
  input \ALUResult_o[1] ;
  input \ALUResult_o[20] ;
  input \ALUResult_o[21] ;
  input \ALUResult_o[22] ;
  input \ALUResult_o[23] ;
  input \ALUResult_o[24] ;
  input \ALUResult_o[25] ;
  input \ALUResult_o[26] ;
  input \ALUResult_o[27] ;
  input \ALUResult_o[28] ;
  input \ALUResult_o[29] ;
  input \ALUResult_o[2] ;
  input \ALUResult_o[30] ;
  input \ALUResult_o[31] ;
  input \ALUResult_o[3] ;
  input \ALUResult_o[4] ;
  input \ALUResult_o[5] ;
  input \ALUResult_o[6] ;
  input \ALUResult_o[7] ;
  input \ALUResult_o[8] ;
  input \ALUResult_o[9] ;
  input \RDData_i[0] ;
  input \RDData_i[10] ;
  input \RDData_i[11] ;
  input \RDData_i[12] ;
  input \RDData_i[13] ;
  input \RDData_i[14] ;
  input \RDData_i[15] ;
  input \RDData_i[16] ;
  input \RDData_i[17] ;
  input \RDData_i[18] ;
  input \RDData_i[19] ;
  input \RDData_i[1] ;
  input \RDData_i[20] ;
  input \RDData_i[21] ;
  input \RDData_i[22] ;
  input \RDData_i[23] ;
  input \RDData_i[24] ;
  input \RDData_i[25] ;
  input \RDData_i[26] ;
  input \RDData_i[27] ;
  input \RDData_i[28] ;
  input \RDData_i[29] ;
  input \RDData_i[2] ;
  input \RDData_i[30] ;
  input \RDData_i[31] ;
  input \RDData_i[3] ;
  input \RDData_i[4] ;
  input \RDData_i[5] ;
  input \RDData_i[6] ;
  input \RDData_i[7] ;
  input \RDData_i[8] ;
  input \RDData_i[9] ;
  input \RDData_o[0] ;
  input \RDData_o[10] ;
  input \RDData_o[11] ;
  input \RDData_o[12] ;
  input \RDData_o[13] ;
  input \RDData_o[14] ;
  input \RDData_o[15] ;
  input \RDData_o[16] ;
  input \RDData_o[17] ;
  input \RDData_o[18] ;
  input \RDData_o[19] ;
  input \RDData_o[1] ;
  input \RDData_o[20] ;
  input \RDData_o[21] ;
  input \RDData_o[22] ;
  input \RDData_o[23] ;
  input \RDData_o[24] ;
  input \RDData_o[25] ;
  input \RDData_o[26] ;
  input \RDData_o[27] ;
  input \RDData_o[28] ;
  input \RDData_o[29] ;
  input \RDData_o[2] ;
  input \RDData_o[30] ;
  input \RDData_o[31] ;
  input \RDData_o[3] ;
  input \RDData_o[4] ;
  input \RDData_o[5] ;
  input \RDData_o[6] ;
  input \RDData_o[7] ;
  input \RDData_o[8] ;
  input \RDData_o[9] ;
  input \RDaddr_i[0] ;
  input \RDaddr_i[1] ;
  input \RDaddr_i[2] ;
  input \RDaddr_i[3] ;
  input \RDaddr_i[4] ;
  input \RDaddr_o[0] ;
  input \RDaddr_o[1] ;
  input \RDaddr_o[2] ;
  input \RDaddr_o[3] ;
  input \RDaddr_o[4] ;
  input \VALUResult_i[0] ;
  input \VALUResult_i[10] ;
  input \VALUResult_i[11] ;
  input \VALUResult_i[12] ;
  input \VALUResult_i[13] ;
  input \VALUResult_i[14] ;
  input \VALUResult_i[15] ;
  input \VALUResult_i[16] ;
  input \VALUResult_i[17] ;
  input \VALUResult_i[18] ;
  input \VALUResult_i[19] ;
  input \VALUResult_i[1] ;
  input \VALUResult_i[20] ;
  input \VALUResult_i[21] ;
  input \VALUResult_i[22] ;
  input \VALUResult_i[23] ;
  input \VALUResult_i[24] ;
  input \VALUResult_i[25] ;
  input \VALUResult_i[26] ;
  input \VALUResult_i[27] ;
  input \VALUResult_i[28] ;
  input \VALUResult_i[29] ;
  input \VALUResult_i[2] ;
  input \VALUResult_i[30] ;
  input \VALUResult_i[31] ;
  input \VALUResult_i[3] ;
  input \VALUResult_i[4] ;
  input \VALUResult_i[5] ;
  input \VALUResult_i[6] ;
  input \VALUResult_i[7] ;
  input \VALUResult_i[8] ;
  input \VALUResult_i[9] ;
  input \VALUResult_o[0] ;
  input \VALUResult_o[10] ;
  input \VALUResult_o[11] ;
  input \VALUResult_o[12] ;
  input \VALUResult_o[13] ;
  input \VALUResult_o[14] ;
  input \VALUResult_o[15] ;
  input \VALUResult_o[16] ;
  input \VALUResult_o[17] ;
  input \VALUResult_o[18] ;
  input \VALUResult_o[19] ;
  input \VALUResult_o[1] ;
  input \VALUResult_o[20] ;
  input \VALUResult_o[21] ;
  input \VALUResult_o[22] ;
  input \VALUResult_o[23] ;
  input \VALUResult_o[24] ;
  input \VALUResult_o[25] ;
  input \VALUResult_o[26] ;
  input \VALUResult_o[27] ;
  input \VALUResult_o[28] ;
  input \VALUResult_o[29] ;
  input \VALUResult_o[2] ;
  input \VALUResult_o[30] ;
  input \VALUResult_o[31] ;
  input \VALUResult_o[3] ;
  input \VALUResult_o[4] ;
  input \VALUResult_o[5] ;
  input \VALUResult_o[6] ;
  input \VALUResult_o[7] ;
  input \VALUResult_o[8] ;
  input \VALUResult_o[9] ;
  input \instr_i[0] ;
  input \instr_i[10] ;
  input \instr_i[11] ;
  input \instr_i[12] ;
  input \instr_i[13] ;
  input \instr_i[14] ;
  input \instr_i[15] ;
  input \instr_i[16] ;
  input \instr_i[17] ;
  input \instr_i[18] ;
  input \instr_i[19] ;
  input \instr_i[1] ;
  input \instr_i[20] ;
  input \instr_i[21] ;
  input \instr_i[22] ;
  input \instr_i[23] ;
  input \instr_i[24] ;
  input \instr_i[25] ;
  input \instr_i[26] ;
  input \instr_i[27] ;
  input \instr_i[28] ;
  input \instr_i[29] ;
  input \instr_i[2] ;
  input \instr_i[30] ;
  input \instr_i[31] ;
  input \instr_i[3] ;
  input \instr_i[4] ;
  input \instr_i[5] ;
  input \instr_i[6] ;
  input \instr_i[7] ;
  input \instr_i[8] ;
  input \instr_i[9] ;
  input \instr_o[0] ;
  input \instr_o[10] ;
  input \instr_o[11] ;
  input \instr_o[12] ;
  input \instr_o[13] ;
  input \instr_o[14] ;
  input \instr_o[15] ;
  input \instr_o[16] ;
  input \instr_o[17] ;
  input \instr_o[18] ;
  input \instr_o[19] ;
  input \instr_o[1] ;
  input \instr_o[20] ;
  input \instr_o[21] ;
  input \instr_o[22] ;
  input \instr_o[23] ;
  input \instr_o[24] ;
  input \instr_o[25] ;
  input \instr_o[26] ;
  input \instr_o[27] ;
  input \instr_o[28] ;
  input \instr_o[29] ;
  input \instr_o[2] ;
  input \instr_o[30] ;
  input \instr_o[31] ;
  input \instr_o[3] ;
  input \instr_o[4] ;
  input \instr_o[5] ;
  input \instr_o[6] ;
  input \instr_o[7] ;
  input \instr_o[8] ;
  input \instr_o[9] ;
  input \pc_i[0] ;
  input \pc_i[10] ;
  input \pc_i[11] ;
  input \pc_i[12] ;
  input \pc_i[13] ;
  input \pc_i[14] ;
  input \pc_i[15] ;
  input \pc_i[16] ;
  input \pc_i[17] ;
  input \pc_i[18] ;
  input \pc_i[19] ;
  input \pc_i[1] ;
  input \pc_i[20] ;
  input \pc_i[21] ;
  input \pc_i[22] ;
  input \pc_i[23] ;
  input \pc_i[24] ;
  input \pc_i[25] ;
  input \pc_i[26] ;
  input \pc_i[27] ;
  input \pc_i[28] ;
  input \pc_i[29] ;
  input \pc_i[2] ;
  input \pc_i[30] ;
  input \pc_i[31] ;
  input \pc_i[3] ;
  input \pc_i[4] ;
  input \pc_i[5] ;
  input \pc_i[6] ;
  input \pc_i[7] ;
  input \pc_i[8] ;
  input \pc_i[9] ;
  input \pc_o[0] ;
  input \pc_o[10] ;
  input \pc_o[11] ;
  input \pc_o[12] ;
  input \pc_o[13] ;
  input \pc_o[14] ;
  input \pc_o[15] ;
  input \pc_o[16] ;
  input \pc_o[17] ;
  input \pc_o[18] ;
  input \pc_o[19] ;
  input \pc_o[1] ;
  input \pc_o[20] ;
  input \pc_o[21] ;
  input \pc_o[22] ;
  input \pc_o[23] ;
  input \pc_o[24] ;
  input \pc_o[25] ;
  input \pc_o[26] ;
  input \pc_o[27] ;
  input \pc_o[28] ;
  input \pc_o[29] ;
  input \pc_o[2] ;
  input \pc_o[30] ;
  input \pc_o[31] ;
  input \pc_o[3] ;
  input \pc_o[4] ;
  input \pc_o[5] ;
  input \pc_o[6] ;
  input \pc_o[7] ;
  input \pc_o[8] ;
  input \pc_o[9] ;
  input clk_i ;
  input start_i ;
  input zero_i ;
  input zero_o ;
  NOT _170_ (
    .A(start_i),
    .Y(_169_)
  );
  NOT _171_ (
    .A(start_i),
    .Y(_000_)
  );
  NOT _172_ (
    .A(start_i),
    .Y(_001_)
  );
  NOT _173_ (
    .A(start_i),
    .Y(_002_)
  );
  NOT _174_ (
    .A(start_i),
    .Y(_003_)
  );
  NOT _175_ (
    .A(start_i),
    .Y(_004_)
  );
  NOT _176_ (
    .A(start_i),
    .Y(_005_)
  );
  NOT _177_ (
    .A(start_i),
    .Y(_006_)
  );
  NOT _178_ (
    .A(start_i),
    .Y(_007_)
  );
  NOT _179_ (
    .A(start_i),
    .Y(_008_)
  );
  NOT _180_ (
    .A(start_i),
    .Y(_009_)
  );
  NOT _181_ (
    .A(start_i),
    .Y(_010_)
  );
  NOT _182_ (
    .A(start_i),
    .Y(_011_)
  );
  NOT _183_ (
    .A(start_i),
    .Y(_012_)
  );
  NOT _184_ (
    .A(start_i),
    .Y(_013_)
  );
  NOT _185_ (
    .A(start_i),
    .Y(_014_)
  );
  NOT _186_ (
    .A(start_i),
    .Y(_015_)
  );
  NOT _187_ (
    .A(start_i),
    .Y(_016_)
  );
  NOT _188_ (
    .A(start_i),
    .Y(_017_)
  );
  NOT _189_ (
    .A(start_i),
    .Y(_018_)
  );
  NOT _190_ (
    .A(start_i),
    .Y(_019_)
  );
  NOT _191_ (
    .A(start_i),
    .Y(_020_)
  );
  NOT _192_ (
    .A(start_i),
    .Y(_021_)
  );
  NOT _193_ (
    .A(start_i),
    .Y(_022_)
  );
  NOT _194_ (
    .A(start_i),
    .Y(_023_)
  );
  NOT _195_ (
    .A(start_i),
    .Y(_024_)
  );
  NOT _196_ (
    .A(start_i),
    .Y(_025_)
  );
  NOT _197_ (
    .A(start_i),
    .Y(_026_)
  );
  NOT _198_ (
    .A(start_i),
    .Y(_027_)
  );
  NOT _199_ (
    .A(start_i),
    .Y(_028_)
  );
  NOT _200_ (
    .A(start_i),
    .Y(_029_)
  );
  NOT _201_ (
    .A(start_i),
    .Y(_030_)
  );
  NOT _202_ (
    .A(start_i),
    .Y(_031_)
  );
  NOT _203_ (
    .A(start_i),
    .Y(_032_)
  );
  NOT _204_ (
    .A(start_i),
    .Y(_033_)
  );
  NOT _205_ (
    .A(start_i),
    .Y(_034_)
  );
  NOT _206_ (
    .A(start_i),
    .Y(_035_)
  );
  NOT _207_ (
    .A(start_i),
    .Y(_036_)
  );
  NOT _208_ (
    .A(start_i),
    .Y(_037_)
  );
  NOT _209_ (
    .A(start_i),
    .Y(_038_)
  );
  NOT _210_ (
    .A(start_i),
    .Y(_039_)
  );
  NOT _211_ (
    .A(start_i),
    .Y(_040_)
  );
  NOT _212_ (
    .A(start_i),
    .Y(_041_)
  );
  NOT _213_ (
    .A(start_i),
    .Y(_042_)
  );
  NOT _214_ (
    .A(start_i),
    .Y(_043_)
  );
  NOT _215_ (
    .A(start_i),
    .Y(_044_)
  );
  NOT _216_ (
    .A(start_i),
    .Y(_045_)
  );
  NOT _217_ (
    .A(start_i),
    .Y(_046_)
  );
  NOT _218_ (
    .A(start_i),
    .Y(_047_)
  );
  NOT _219_ (
    .A(start_i),
    .Y(_048_)
  );
  NOT _220_ (
    .A(start_i),
    .Y(_049_)
  );
  NOT _221_ (
    .A(start_i),
    .Y(_050_)
  );
  NOT _222_ (
    .A(start_i),
    .Y(_051_)
  );
  NOT _223_ (
    .A(start_i),
    .Y(_052_)
  );
  NOT _224_ (
    .A(start_i),
    .Y(_053_)
  );
  NOT _225_ (
    .A(start_i),
    .Y(_054_)
  );
  NOT _226_ (
    .A(start_i),
    .Y(_055_)
  );
  NOT _227_ (
    .A(start_i),
    .Y(_056_)
  );
  NOT _228_ (
    .A(start_i),
    .Y(_057_)
  );
  NOT _229_ (
    .A(start_i),
    .Y(_058_)
  );
  NOT _230_ (
    .A(start_i),
    .Y(_059_)
  );
  NOT _231_ (
    .A(start_i),
    .Y(_060_)
  );
  NOT _232_ (
    .A(start_i),
    .Y(_061_)
  );
  NOT _233_ (
    .A(start_i),
    .Y(_062_)
  );
  NOT _234_ (
    .A(start_i),
    .Y(_063_)
  );
  NOT _235_ (
    .A(start_i),
    .Y(_064_)
  );
  NOT _236_ (
    .A(start_i),
    .Y(_065_)
  );
  NOT _237_ (
    .A(start_i),
    .Y(_066_)
  );
  NOT _238_ (
    .A(start_i),
    .Y(_067_)
  );
  NOT _239_ (
    .A(start_i),
    .Y(_068_)
  );
  NOT _240_ (
    .A(start_i),
    .Y(_069_)
  );
  NOT _241_ (
    .A(start_i),
    .Y(_070_)
  );
  NOT _242_ (
    .A(start_i),
    .Y(_071_)
  );
  NOT _243_ (
    .A(start_i),
    .Y(_072_)
  );
  NOT _244_ (
    .A(start_i),
    .Y(_073_)
  );
  NOT _245_ (
    .A(start_i),
    .Y(_074_)
  );
  NOT _246_ (
    .A(start_i),
    .Y(_075_)
  );
  NOT _247_ (
    .A(start_i),
    .Y(_076_)
  );
  NOT _248_ (
    .A(start_i),
    .Y(_077_)
  );
  NOT _249_ (
    .A(start_i),
    .Y(_078_)
  );
  NOT _250_ (
    .A(start_i),
    .Y(_079_)
  );
  NOT _251_ (
    .A(start_i),
    .Y(_080_)
  );
  NOT _252_ (
    .A(start_i),
    .Y(_081_)
  );
  NOT _253_ (
    .A(start_i),
    .Y(_082_)
  );
  NOT _254_ (
    .A(start_i),
    .Y(_083_)
  );
  NOT _255_ (
    .A(start_i),
    .Y(_084_)
  );
  NOT _256_ (
    .A(start_i),
    .Y(_085_)
  );
  NOT _257_ (
    .A(start_i),
    .Y(_086_)
  );
  NOT _258_ (
    .A(start_i),
    .Y(_087_)
  );
  NOT _259_ (
    .A(start_i),
    .Y(_088_)
  );
  NOT _260_ (
    .A(start_i),
    .Y(_089_)
  );
  NOT _261_ (
    .A(start_i),
    .Y(_090_)
  );
  NOT _262_ (
    .A(start_i),
    .Y(_091_)
  );
  NOT _263_ (
    .A(start_i),
    .Y(_092_)
  );
  NOT _264_ (
    .A(start_i),
    .Y(_093_)
  );
  NOT _265_ (
    .A(start_i),
    .Y(_094_)
  );
  NOT _266_ (
    .A(start_i),
    .Y(_095_)
  );
  NOT _267_ (
    .A(start_i),
    .Y(_096_)
  );
  NOT _268_ (
    .A(start_i),
    .Y(_097_)
  );
  NOT _269_ (
    .A(start_i),
    .Y(_098_)
  );
  NOT _270_ (
    .A(start_i),
    .Y(_099_)
  );
  NOT _271_ (
    .A(start_i),
    .Y(_100_)
  );
  NOT _272_ (
    .A(start_i),
    .Y(_101_)
  );
  NOT _273_ (
    .A(start_i),
    .Y(_102_)
  );
  NOT _274_ (
    .A(start_i),
    .Y(_103_)
  );
  NOT _275_ (
    .A(start_i),
    .Y(_104_)
  );
  NOT _276_ (
    .A(start_i),
    .Y(_105_)
  );
  NOT _277_ (
    .A(start_i),
    .Y(_106_)
  );
  NOT _278_ (
    .A(start_i),
    .Y(_107_)
  );
  NOT _279_ (
    .A(start_i),
    .Y(_108_)
  );
  NOT _280_ (
    .A(start_i),
    .Y(_109_)
  );
  NOT _281_ (
    .A(start_i),
    .Y(_110_)
  );
  NOT _282_ (
    .A(start_i),
    .Y(_111_)
  );
  NOT _283_ (
    .A(start_i),
    .Y(_112_)
  );
  NOT _284_ (
    .A(start_i),
    .Y(_113_)
  );
  NOT _285_ (
    .A(start_i),
    .Y(_114_)
  );
  NOT _286_ (
    .A(start_i),
    .Y(_115_)
  );
  NOT _287_ (
    .A(start_i),
    .Y(_116_)
  );
  NOT _288_ (
    .A(start_i),
    .Y(_117_)
  );
  NOT _289_ (
    .A(start_i),
    .Y(_118_)
  );
  NOT _290_ (
    .A(start_i),
    .Y(_119_)
  );
  NOT _291_ (
    .A(start_i),
    .Y(_120_)
  );
  NOT _292_ (
    .A(start_i),
    .Y(_121_)
  );
  NOT _293_ (
    .A(start_i),
    .Y(_122_)
  );
  NOT _294_ (
    .A(start_i),
    .Y(_123_)
  );
  NOT _295_ (
    .A(start_i),
    .Y(_124_)
  );
  NOT _296_ (
    .A(start_i),
    .Y(_125_)
  );
  NOT _297_ (
    .A(start_i),
    .Y(_126_)
  );
  NOT _298_ (
    .A(start_i),
    .Y(_127_)
  );
  NOT _299_ (
    .A(start_i),
    .Y(_128_)
  );
  NOT _300_ (
    .A(start_i),
    .Y(_129_)
  );
  NOT _301_ (
    .A(start_i),
    .Y(_130_)
  );
  NOT _302_ (
    .A(start_i),
    .Y(_131_)
  );
  NOT _303_ (
    .A(start_i),
    .Y(_132_)
  );
  NOT _304_ (
    .A(start_i),
    .Y(_133_)
  );
  NOT _305_ (
    .A(start_i),
    .Y(_134_)
  );
  NOT _306_ (
    .A(start_i),
    .Y(_135_)
  );
  NOT _307_ (
    .A(start_i),
    .Y(_136_)
  );
  NOT _308_ (
    .A(start_i),
    .Y(_137_)
  );
  NOT _309_ (
    .A(start_i),
    .Y(_138_)
  );
  NOT _310_ (
    .A(start_i),
    .Y(_139_)
  );
  NOT _311_ (
    .A(start_i),
    .Y(_140_)
  );
  NOT _312_ (
    .A(start_i),
    .Y(_141_)
  );
  NOT _313_ (
    .A(start_i),
    .Y(_142_)
  );
  NOT _314_ (
    .A(start_i),
    .Y(_143_)
  );
  NOT _315_ (
    .A(start_i),
    .Y(_144_)
  );
  NOT _316_ (
    .A(start_i),
    .Y(_145_)
  );
  NOT _317_ (
    .A(start_i),
    .Y(_146_)
  );
  NOT _318_ (
    .A(start_i),
    .Y(_147_)
  );
  NOT _319_ (
    .A(start_i),
    .Y(_148_)
  );
  NOT _320_ (
    .A(start_i),
    .Y(_149_)
  );
  NOT _321_ (
    .A(start_i),
    .Y(_150_)
  );
  NOT _322_ (
    .A(start_i),
    .Y(_151_)
  );
  NOT _323_ (
    .A(start_i),
    .Y(_152_)
  );
  NOT _324_ (
    .A(start_i),
    .Y(_153_)
  );
  NOT _325_ (
    .A(start_i),
    .Y(_154_)
  );
  NOT _326_ (
    .A(start_i),
    .Y(_155_)
  );
  NOT _327_ (
    .A(start_i),
    .Y(_156_)
  );
  NOT _328_ (
    .A(start_i),
    .Y(_157_)
  );
  NOT _329_ (
    .A(start_i),
    .Y(_158_)
  );
  NOT _330_ (
    .A(start_i),
    .Y(_159_)
  );
  NOT _331_ (
    .A(start_i),
    .Y(_160_)
  );
  NOT _332_ (
    .A(start_i),
    .Y(_161_)
  );
  NOT _333_ (
    .A(start_i),
    .Y(_162_)
  );
  NOT _334_ (
    .A(start_i),
    .Y(_163_)
  );
  NOT _335_ (
    .A(start_i),
    .Y(_164_)
  );
  NOT _336_ (
    .A(start_i),
    .Y(_165_)
  );
  NOT _337_ (
    .A(start_i),
    .Y(_166_)
  );
  NOT _338_ (
    .A(start_i),
    .Y(_167_)
  );
  NOT _339_ (
    .A(start_i),
    .Y(_168_)
  );
endmodule
